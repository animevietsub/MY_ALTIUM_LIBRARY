.SUBCKT IIND_COUPLED_4 P11 P12 P21 P22 P31 P32 P41 P42 PARAMS: L1=1u L2=1u L3=1u L4=1u KA=0.98
LL1 P11 P12 {L1}
LL2 P21 P22 {L2}
LL3 P31 P32 {L3}
LL4 P41 P42 {L4}
KKA LL1 LL2 LL3 LL4 {KA}
.ENDS

.SUBCKT IIND_COUPLED_2 P11 P12 P21 P22 PARAMS: L1=1u L2=1u KA=0.98
LL1 P11 P12 {L1}
LL2 P21 P22 {L2}
KKA LL1 LL2 {KA}
.ENDS
