* MCR100-3  SCR  A G K  MCE  7-17-95
*MCE MCR100-3 100V  800mA  pkg:TO-226AA
.SUBCKT MCR100-3 1 2 3
QP  6 4 1  POUT OFF
QN  4 6 5  NOUT OFF
RF  6 4    20MEG
RR  1 4    13.3MEG
RGK 6 5    6.25K
RG  2 6    9.17
RK  3 5    81.3M
DF  6 4    ZF
DR  1 4    ZR
DGK 6 5    ZGK
.MODEL ZF   D (IS=.32F IBV=1U BV=100 RS=3MEG)
.MODEL ZR   D (IS=.32F IBV=1U BV=133)
.MODEL ZGK  D (IS=.32F IBV=1U BV=5)
.MODEL POUT PNP (IS=320F BF=1 CJE=67P)
.MODEL NOUT NPN (IS=320F BF=100 RC=.325
+ CJE=67P CJC=13.4P TF=56.6N TR=8.06U)
.ENDS XMCR1003

* MCR100-4  SCR  A G K  MCE  7-17-95
*MCE MCR100-4 200V  800mA  pkg:TO-226AA
.SUBCKT MCR100-4 1 2 3
QP  6 4 1  POUT OFF
QN  4 6 5  NOUT OFF
RF  6 4    40MEG
RR  1 4    26.6MEG
RGK 6 5    6.25K
RG  2 6    9.17
RK  3 5    81.3M
DF  6 4    ZF
DR  1 4    ZR
DGK 6 5    ZGK
.MODEL ZF   D (IS=.32F IBV=1U BV=200 RS=6MEG)
.MODEL ZR   D (IS=.32F IBV=1U BV=266)
.MODEL ZGK  D (IS=.32F IBV=1U BV=5)
.MODEL POUT PNP (IS=320F BF=1 CJE=67P)
.MODEL NOUT NPN (IS=320F BF=100 RC=.325
+ CJE=67P CJC=13.4P TF=56.6N TR=8.06U)
.ENDS XMCR1004

* MCR100-6  SCR  A G K  MCE  7-17-95
*MCE MCR100-6 400V  800mA  pkg:TO-226AA
.SUBCKT MCR100-6 1 2 3
QP  6 4 1  POUT OFF
QN  4 6 5  NOUT OFF
RF  6 4    80MEG
RR  1 4    53.3MEG
RGK 6 5    6.25K
RG  2 6    9.17
RK  3 5    81.3M
DF  6 4    ZF
DR  1 4    ZR
DGK 6 5    ZGK
.MODEL ZF   D (IS=.32F IBV=1U BV=400 RS=12MEG)
.MODEL ZR   D (IS=.32F IBV=1U BV=533)
.MODEL ZGK  D (IS=.32F IBV=1U BV=5)
.MODEL POUT PNP (IS=320F BF=1 CJE=67P)
.MODEL NOUT NPN (IS=320F BF=100 RC=.325
+ CJE=67P CJC=13.4P TF=56.6N TR=8.06U)
.ENDS XMCR1006

* MCR100-8  SCR  A G K  MCE  7-17-95
*MCE MCR100-8 600V  800mA  pkg:TO-226AA
.SUBCKT MCR100-8 1 2 3
*    TERMINALS:  A G K
*  600 Volt  .8 Amp  SCR  07-17-1995
QP  6 4 1  POUT OFF
QN  4 6 5  NOUT OFF
RF  6 4    120MEG
RR  1 4    80MEG
RGK 6 5    6.25K
RG  2 6    9.17
RK  3 5    81.3M
DF  6 4    ZF
DR  1 4    ZR
DGK 6 5    ZGK
.MODEL ZF   D (IS=.32F IBV=1U BV=600 RS=18MEG)
.MODEL ZR   D (IS=.32F IBV=1U BV=800)
.MODEL ZGK  D (IS=.32F IBV=1U BV=5)
.MODEL POUT PNP (IS=320F BF=1 CJE=67P)
.MODEL NOUT NPN (IS=320F BF=100 RC=.325
+ CJE=67P CJC=13.4P TF=56.6N TR=8.06U)
.ENDS XMCR1008
