*$
**************** Power Discrete MOSFET Electrical Circuit Model *****************
** Product Name: FQD19N10LTM
** N-Channel QFET MOSFET 100V, 15.6A, 100mohm
** Model Type: BSIM3V3
**-------------------------------------------------------------------------------
.SUBCKT FQD19N10L 2 1 3    
*Nom Temp=25 deg C
Dbody 7 5    DbodyMOD
Dbreak 5 11  DbreakMOD
Ebreak 11 7 17 7 110
Lgate 1 9    1.125e-9
Ldrain 2 5   0.966e-10
Lsource 3 7  0.966e-10
RLgate 1 9   11.25
RLdrain 2 5  9.66
RLsource 3 7 9.66
Rgate 9 6    0.5
It 7 17      1
Rbreak 17 7  RbreakMOD 1
.MODEL RbreakMOD RES (TC1=9.28e-4 TC2=-1.03e-6)
.MODEL DbodyMOD D (IS=1.15e-12   N=1.0    RS=1.76e-2  TRS1=1.05e-3  TRS2=1.2e-7 
+ CJO=1.14e-9      M=0.58       VJ=0.46  TT=6.27e-8  XTI=3         EG=1.18)
.MODEL DbreakMOD D (RS=100e-3 TRS1=1.0e-3 TRS2=1e-6)
Rdrain 5 16 RdrainMOD 0.067
.MODEL RdrainMOD RES (TC1=6.02e-3 TC2=1.05e-5)
M_BSIM3 16 6 7 7 Bsim3 W=0.85 L=2.0e-6 NRS=1
.MODEL Bsim3 NMOS (LEVEL=7 VERSION=3.1 MOBMOD=3 CAPMOD=2 PARAMCHK=1 NQSMOD=0
+ TOX=500e-10     XJ=1.4e-6      NCH=1.3e17      
+ U0=700          VSAT=1.0e5     DROUT=1.0     
+ DELTA=0.1       PSCBE2=0       RSH=3.59e-3    
+ VTH0=1.65       VOFF=-0.1      NFACTOR=1.1
+ LINT=3.25e-7    DLC=3.25e-7    FC=0.5
+ CGSO=1.00e-15   CGSL=0         CGDO=2.05e-14 
+ CGDL=1.28e-9    CJ=0           CF=0
+ CKAPPA=0.2      KT1=-1.45      KT2=0
+ UA1=3.8e-9      NJ=10)
.ENDS
*$
********************* Power Discrete MOSFET Thermal Model **********************
** Package: D-PAK
**------------------------------------------------------------------------------
.SUBCKT FQD19N10L_Thermal TH TL
CTHERM1 TH 6 1.01e-5
CTHERM2 6 5  1.25e-3
CTHERM3 5 4  4.52e-3
CTHERM4 4 3  1.85e-2
CTHERM5 3 2  2.40e-2
CTHERM6 2 TL 1.24e-1 
RTHERM1 TH 6 1.76e-2
RTHERM2 6 5  6.06e-2
RTHERM3 5 4  8.90e-2
RTHERM4 4 3  1.83e-1
RTHERM5 3 2  6.200e-1
RTHERM6 2 TL 1.53e+0
.ENDS FQD19N10L_Thermal 
**------------------------------------------------------------------------------
** Creation: Aug.-22-2017   Rev.: 1.0
** ON Semiconductor
*$

