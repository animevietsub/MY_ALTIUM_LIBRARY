* Copyright � Linear Technology Corp. 1998, 1999, 2000.  All rights reserved.
*
.subckt PC817 1 2 3 4
R1 N003 2 2
D1 1 N003 LD
G1 3 N004 N003 2 0.03
C1 1 2 18p
Q1 4 N004 3 NP
.model LD D(Is=1e-20 Cjo=18p Vj=1.2)
.model NP NPN(Bf=100 Vaf=140 Ikf=100m Rc=1 Cjc=19p Cje=7p Cjs=7p)
.ends PC817

