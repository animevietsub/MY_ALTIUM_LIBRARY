* Library of Opamp, Voltage Comparator, Voltage Regulator, Voltage
* Reference Models
*
*  Copyright OrCAD, Inc. 1998 All Rights Reserved.

* $Revision:   1.4  $
* $Author:   rperez  $
* $Date:   28 Oct 1998 13:20:42  $
*
* ---------------------------------------------------------------------------
*** Operational amplifiers

* The parameters in the opamp library were derived from the data sheets for
* each part.  The macromodel used is similar to the one described in:
*
*       Macromodeling of Integrated Circuit Operational Amplifiers
*         by Graeme Boyle, Barry Cohn, Donald Pederson, and James Solomon
*       IEEE Journal of SoliE-State Circuits, Vol. SC-9, no. 6, Dec. 1974
*
* Differences from the reference (above) occur in the output limiting stage
* which was modified to reduce internally generated currents associated with
* output voltage limiting, as well as short-circuit current limiting.
*
* The opamps are modelled at room temperature and do not track changes with
* temperature.  This library file contains models for nominal, not worst case,
* devices.
*$
*-----------------------------------------------------------------------------
*
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt ad648a   1 2 3 4 5
*
  c1   11 12 11.66E-12
  c2    6  7 25.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 127.3E9 -1E3 1E3 130E9 -130E9
  ga    6  0 11 12 157.1E-6
  gcm   0  6 10 99 24.93E-9
  iss  10  4 dc 45.00E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   3 11 6.366E3
  rd2   3 12 6.366E3
  ro1   8  5 50.00E-3
  ro2   7 99 50.00E-3
  rp    3  4 176.5E3
  rss  10 99 4.444E6
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 15
  vln   0 92 dc 15
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=2.500E-12 Beta=548.3E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt AD648B   1 2 3 4 5
*
  c1   11 12 11.66E-12
  c2    6  7 25.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 127.3E9 -1E3 1E3 130E9 -130E9
  ga    6  0 11 12 157.1E-6
  gcm   0  6 10 99 12.47E-9
  iss  10  4 dc 45.00E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   3 11 6.366E3
  rd2   3 12 6.366E3
  ro1   8  5 50.00E-3
  ro2   7 99 50.00E-3
  rp    3  4 176.5E3
  rss  10 99 4.444E6
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 15
  vln   0 92 dc 15
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=1.500E-12 Beta=548.3E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt AD648C   1 2 3 4 5
*
  c1   11 12 11.66E-12
  c2    6  7 25.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 127.3E9 -1E3 1E3 130E9 -130E9
  ga    6  0 11 12 157.1E-6
  gcm   0  6 10 99 7.854E-9
  iss  10  4 dc 45.00E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   3 11 6.366E3
  rd2   3 12 6.366E3
  ro1   8  5 50.00E-3
  ro2   7 99 50.00E-3
  rp    3  4 176.5E3
  rss  10 99 4.444E6
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 15
  vln   0 92 dc 15
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=1.500E-12 Beta=548.3E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt ad741    1 2 3 4 5
*
  c1   11 12 2.645E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 16.32E6 -1E3 1E3 16E6 -16E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.837E3
  re2  14 10 1.837E3
  ree  10 99 13.19E6
  ro1   8  5 45
  ro2   7 99 65
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
*$
*
* MANUFACTURERS PART NO. = HA2-2600-8  (HARRIS)
* SUBTYPE:OP_AMP
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT MODEL OF THE HA2-
* 2600.
* THIS MODEL INCLUDES PARAMETERS WHICH THE MICROSIM-BOYLE MODEL DID NOT.
*
* IT MODELS POWER-UP, POWER-DOWN, AND POWER OFF CONDITIONS,
* SINGLE SUPPLY APPLICATIONS, AC PSRR, DC PSRR, AC CMRR, VSAT, IIB, IIO,
* VIO, ISC, SR, PM, GBP, ICC, AND RO(AC).
*-----------------------------------------------------------------------------
* THE FOLLOWING SPECIFICATIONS ARE SIMULATED IN THE MODEL FOR +/-15 V
* SUPPLIES:
*  VIO = 0.85 MV, VSAT = +13 V, VSAT- = -14 V, IB+ = 2 NA, IB- = -1.3 NA,
*  GBP = 12.4MHZ, PM = 46 DEG, CMRR = 107 DB, RO(AC) = 39 OHMS, ISC+ = 3 MA
*  ISC- = -28 MA, SR+ = 7.5 V/US, SR- = -6.4 V/US
*
* MODIFIED SPECS:
* DC PSRR = 100 DB, AC PSRR MODELED; ISUPPLY = IBIAS + ILOAD, VSAT VARIES WITH
* SUPPLY VOLTAGES, ALSO MODELS SINGLE SUPPLY APPLICATIONS; E.G. VCC+ = 5 V,
* VCC- = 0 V, VSAT+ = 3 V, VSAT- = 5 MV; POWER NOT CONNECTED MODELED; POWER-
* UP  AND POWER-DOWN MODELED. INPUT BIAS CURRENT CAN BE + OR -.
*
* THIS MODEL CAN BE USED WITH A .TEMP CARD OVER THE TEMPERATURE RANGE
* OF  -55 C TO 125 C.
*
* THE FOLLOWING PARAMETERS ARE INSENSITIVE TO TEMPERATURE CHANGES AND
* ARE  SIMULATED ACCURATELY BY THE MODEL: CMRR  GAIN  ICC  PSRR  SR
* OVERDRIVE  RECOVERY TIME   OUTPUT VOLTAGE SWING  IIB  IIO
*
* THE FOLLOWING PARAMETERS ARE TEMPERATURE DEPENDENT AND ARE
* SIMULATED BY THE MODEL:  ISC  VIO
*
*
* CONNECTIONS:    NON-INVERTING INPUT
*                 | INVERTING INPUT
*                 | | POSITIVE POWER SUPPLY
*                 | | | NEGATIVE POWER SUPPLY
*                 | | |  | OUTPUT
*                 | | |  |   |  GND(REFERENCE)
*                 | | |  |   |   |
.SUBCKT HA-2600   1 2 3A 4A  5  100
*
* DC PSRR FIX
Q1 11 16 13 HA2600QA
EPSRR- 16 2 TABLE {-V(4)} = (0,150U) (20,-50U)
Q2 12 15 14 HA2600QB
EPSRR+ 1 15 TABLE {V(3)} = (0,150U) (20,-50U)
*
*INPUT CURRENT COMPENSATION
IBX1 100 16 6.3N
IBX2 100 15 2.99N
*
RC1 3 11 1276
RC2 3 12 1276
C1 11 12 6.6519P
RE1 13 10 573
RE2 14 10 573
GIEE 10 4 TABLE {V(3,4)} = (0,0) (2,0) (3,73.6U)
CE 10 100 1.464P
RE 10 100 2.717MEG
RP 3 4 9913
*
* CMRR FIX
GCM1 100 83 10 100 1
RCM1 83 84 1
LCM1 84 100 1.592U
GCM2 100 85 83 100 1
RCM2 85 86 1
LCM2 86 100 0.1592U
RCM3 86 100 10
GCM 100 21 85 100 3.5N
*
GA 21 100 11 12 783.7U
*
* PSRR VS FREQ FIX
GPSRR- 21 100 88 100 1
GVP- 100 88 4 100 1
RVP- 88 100 1
LVP- 88 100 10P
GPSRR+ 21 100 89 100 1
GVP+ 100 89 3 100 1
RVP+ 89 100 1
LVP+ 89 100 0.1P
*
R2 21 100 100K
C2 21 22 10P
GB 22 100 21 100 1359
RO2 22 100 41
D1 22 31 HA2600DA
D2 31 22 HA2600DC
EC 31 100 5 100 1.0
*
* I(VCC) FIX
RO1 22 6 39
VIOUT 6 5 0
D5 3 7 HA2600DB
R5 7 100 1MEG
F5 7 100 VIOUT 1
D6 8 4 HA2600DB
R6 8 100 1MEG
F6 8 100 VIOUT 1
*
* POWER OFF FIX
VIVP+ 3A 3
WVP+ 3 3B VIVP+ CL1
VIVP- 4 4A
WVP- 4 4B VIVP- CL1
.MODEL CL1 ISWITCH(
+        RON = 0.1
+       ROFF = 10MEG
+        ION = 0.5U
+       IOFF = 1N
+ )
*
* CLIPPING FIX
D3 5 24 HA2600DB
EVC 3B 24 TABLE {V(3)} = (0,0.81089) (5,2.81089)
D4 25 5 HA2600DB
EVE 25 4B TABLE {-V(4)} = (0,0.80648) (5,1.80648)
*
.MODEL HA2600DA D (
+         IS = 1.8E-18
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL HA2600DC D (
+         IS = 4.581F
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL HA2600DB D (
+         IS = 0.8F
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL HA2600QA NPN (
+         IS = 0.827F
+         BF = 7360
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
.MODEL HA2600QB NPN (
+         IS = 0.8F
+         BF = 7360
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
.ENDS HA-2600
*$
*
* MANUFACTURERS PART NO. = HA7-2720-8  (HARRIS)
* SUBTYPE: OP_AMP
* THIS FILE CONTAINS 1 PRE-RAD MODEL AT 27 C OF THE HA7-2720.
*
*
* THIS MACROMODEL IS DERIVED FROM A MODIFIED BOYLE MACROMODEL STRUCTURE.
*
* PARAMETERS THAT VARY WITH ISET INCLUDE: GAIN BANDWIDTH PRODUCT; POWER
* DISSIPATED; CMRR; SHORT CIRCUIT CURRENT; SLEW RATE; OUTPUT RESISTANCE
*
.SUBCKT HA-2720   1   2   3   4   5   27   100
*              +IN   |   |   |   |   |     |
*                  -IN   |   |   |   |     |
*                      +VCC  |   |   |     |
*                          -VCC  |   |     |
*                               OUT  |     |
*                                  ISET    |
*                                       GND(REFERENCE)
C1 11 12 0.8P
C2 6 7 10P
DC 5 53 DX
DE 54 5 DX
DLP 90 91 DX
DLN 92 90 DX
DP 4 3 DX
EGND 99 100 POLY(2) (3,100) (4,100) 0 0.5 0.5
FB 7 99 POLY(5) VB VC VE VLP VLN 0 1.061E9 -9E8 1E9 1E9 -1E9
GA 6 100 11 12 9.425U
GCM 100 6 10 99 298P
FIEE 10 4 VSET 0.667
HLIM 90 100 VLIM 10K
Q1 11 2 13 QX
Q2 12 1 14 QX
R2 6 9 10K
RC1 3 11 106.1K
RC2 3 12 106.1K
RE1 13 10 54.4K
RE2 14 10 54.4K
REE 10 99 200MEG
RO1  8 5 10
RO2  7 99 10
VB 9 100 DC 0
VC 3 53 DC 1
VE 54 4 DC 1
VLIM 7 8  DC 0
VLP 91 89 DC 0
VLN 88 92 DC 0
*
* ADDITIONAL MODEL COMPONENTS
*
D1 3 25 DX
D2 25 26 DX
VSET 26 27 DC 0
FDISP 3 4 VSET 13
HLP 89 100 VSET 3.33MEG
HLN 100 88 VSET 3.33MEG
*
.MODEL DX D(
+         IS = 800E-18
+         RS = 1
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.MODEL QX NPN(
+         IS = 800E-18
+         BF = 250
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.ENDS HA-2720
*$
*
* MANUFACTURERS PART NO. = HA5154/883  (HARRIS)
* SUBTYPE: OP_AMP
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT MODEL OF THE HA5154.
*
* IT MODELS POWER-UP, POWER-DOWN, AND POWER OFF CONDITIONS,
* SINGLE SUPPLY APPLICATIONS, AC PSRR, DC PSRR, AC CMRR, VSAT, IIB, IIO,
* VIO, ISC, SR, PM, GBP, ICC, AND RO(AC).
*----------------------------------------------------------------------------
* THE FOLLOWING SPECIFICATIONS ARE SIMULATED IN THE MODEL FOR +/-15 V
* SUPPLIES:
*  VIO = 0.4 MV, VSAT = +13.5 V, VSAT- = -13.8 V,IB+ = 113.5 NA,IB- = -111.6NA
*  GBP = 1.26MHZ, PM = 78 DEG, CMRR = 102 DB, RO(AC) = 317 OHMS, ISC+ = 8.8 MA
*  ISC- = -3.4 MA, SR+ = 6.66 V/US, SR- = -7.4 V/US
*
* MODIFIED SPECS:
* DC PSRR = 100 DB, AC PSRR MODELED; ISUPPLY = IBIAS + ILOAD, VSAT VARIES WITH
* SUPPLY VOLTAGES, ALSO MODELS SINGLE SUPPLY APPLICATIONS; E.G. VCC+ = 5 V,
* VCC- = 0 V, VSAT+ = 3 V, VSAT- = 5 MV; POWER NOT CONNECTED MODELED; POWER-
* UP  AND POWER-DOWN MODELED. INPUT BIAS CURRENT CAN BE + OR -.
*
* THIS MODEL CAN BE USED WITH A .TEMP CARD OVER THE TEMPERATURE RANGE
* OF  -55 C TO 125 C.
*
* THE FOLLOWING PARAMETERS ARE INSENSITIVE TO TEMPERATURE CHANGES AND
* ARE  SIMULATED ACCURATELY BY THE MODEL: CMRR  GAIN  ICC  PSRR  SR
* OVERDRIVE  RECOVERY TIME   OUTPUT VOLTAGE SWING  IIB  IIO
*
* THE FOLLOWING PARAMETERS ARE TEMPERATURE DEPENDENT AND ARE
* SIMULATED  BY THE MODEL:  ISC  VIO
*
*
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | |  | OUTPUT
*                | | |  |   |   GND(REFERENCE)
*                | | |  |   |    |
.SUBCKT HA-5154   1 2 3A 4A  5A  100
*
* DC PSRR FIX
Q1 11 16 13 HA5154QA
EPSRR- 16 2 TABLE {-V(4)} = (0,150U) (20,-50U)
Q2 12 15 14 HA5154QB
EPSRR+ 1 15 TABLE {V(3)} = (0,150U) (20,-50U)
*
*INPUT CURRENT COMPENSATION
IBX1 16 100 186N
IBX2 15 100 188N
*
RC1 4 11 12.25K
RC2 4 12 12.25K
C1 11 12 1.072P
RE1 13 10 11.56K
RE2 14 10 11.56K
GIEE 3 10 TABLE {V(3,4)} = (0,0) (2,0) (3,75U)
CE 10 100 0.838P
RE 10 100 2.67MEG
*
* SUPPLY CURRENT FOR 1/4 CURRENT OF IC.
* PLACE AN RP IN PARALLEL FOR EACH UNUSED OPAMP ON IC.
*
RP 3 4 171K
*
* CMRR FIX
GCM1 100 83 10 100 1
RCM1 83 84 1
LCM1 84 100 15.92U
GCM2 100 85 83 100 1
RCM2 85 86 1
LCM2 86 100 1.592U
RCM3 86 100 10
GCM 100 21 85 100 0.648N
*
GA 21 100 11 12 81.63U
*
* PSRR VS FREQ FIX
GPSRR- 21 100 88 100 1
GVP- 100 88 4 100 1
RVP- 88 100 1
LVP- 88 100 0.10P
GPSRR+ 21 100 89 100 1
GVP+ 100 89 3 100 1
RVP+ 89 100 1
LVP+ 89 100 10P
*
R2 21 100 100K
C2 21 22 10P
GB 22 100 21 100 297.89
RO2 22 100 83
D1 22 31 HA5154DA
D2 31 22 HA5154DC
EC 31 100 5 100 1.0
*
* I(VCC) FIX
RO1 22 6 217
VIOUT 6 5 0
D5 3 7 HA5154DB
R5 7 100 1MEG
F5 7 100 VIOUT 1
D6 8 4 HA5154DB
R6 8 100 1MEG
F6 8 100 VIOUT 1
*
*EXTERNAL RO AT VO
RO3 5 5A 100
*
* POWER OFF FIX
VIVP+ 3A 3
WVP+ 3 3B VIVP+ CL1
VIVP- 4 4A
WVP- 4 4B VIVP- CL1
.MODEL CL1 ISWITCH(
+        RON = 0.1
+       ROFF = 50MEG
+        ION = 0.5U
+       IOFF = 1N
+ )
*
* CLIPPING FIX
D3 5 24 HA5154DB
EVC 3B 24 TABLE {V(3)} = (0,0.77655) (3,2.17655)
D4 25 5 HA5154DB
EVE 25 4B TABLE {-V(4)} = (0,0.751956) (3,1.751956)
*
.MODEL HA5154DA D (
+         IS = 19.02E-30
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL HA5154DC D (
+         IS = 908.77P
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL HA5154DB D (
+         IS = 0.8F
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL HA5154QA NPN (
+         IS = 0.7879F
+         BF = 500
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
.MODEL HA5154QB NPN (
+         IS = 0.8F
+         BF = 500
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
.ENDS HA-5154
*$
*
* MANUFACTURERS PART NO. = HS3516RH  (HARRIS)
* SUBTYPE:OP_AMP
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT MODEL OF THE HS3516.
*
* IT MODELS POWER-UP, POWER-DOWN, AND POWER OFF CONDITIONS,
* SINGLE SUPPLY APPLICATIONS, AC PSRR, DC PSRR, AC CMRR, VSAT, IIB, IIO,
* VIO, ISC, SR, PM, GBP, ICC, AND RO(AC). THE VOLTAGE CLAMPING PIN HAS
* BEEN MODELED. IT HAS BEEN COMMENTED OUT WITH THE * SYMBOL BECAUSE IT
* CAN  CAUSE CONVERGENCE PROBLEMS. TO ADD TO THE MODEL ADD PIN 9 ON THE
*.SUBCKT  LINE AND REMOVE THE * FROM THE LINES DEFINING THE CLAMP PIN IN THE
* MODEL.  IF IT CAUSES A CONVERGENCE PROBLEM USE ITL4=300 IN THE .OPTION
* STATEMENT.
*-----------------------------------------------------------------------------
* THE FOLLOWING SPECIFICATIONS ARE SIMULATED IN THE MODEL FOR +/-15 V
* SUPPLIES:
*  VIO = 0.52 MV, VSAT = +13.5 V, VSAT- = -12.6 V, IB = 14.8 NA, IIO = -6 NA
*  GBP = 11MHZ, PM = 47 DEG, CMRR = 107 DB, RO(AC) = 30 OHMS, ISC+ = 26 MA
*  ISC- = -27 MA, SR+ = 23.4 V/US, SR- = -21 V/US
*
* MODIFIED SPECS:
* DC PSRR = 100 DB, AC PSRR MODELED; ISUPPLY = IBIAS + ILOAD, VSAT VARIES WITH
* SUPPLY VOLTAGES, ALSO MODELS SINGLE SUPPLY APPLICATIONS; E.G. VCC+ = 5 V,
* VCC- = 0 V, VSAT+ = 3 V, VSAT- = 5 MV; POWER NOT CONNECTED MODELED; POWER-
* UP  AND POWER-DOWN MODELED.
*
* THIS MODEL CAN BE USED WITH A .TEMP CARD OVER THE TEMPERATURE RANGE
* OF  -55 C TO 125 C.
*
* THE FOLLOWING PARAMETERS ARE INSENSITIVE TO TEMPERATURE CHANGES AND
* ARE  SIMULATED ACCURATELY BY THE MODEL: CMRR  GAIN  ICC  PSRR  SR
* OVERDRIVE  RECOVERY TIME   OUTPUT VOLTAGE SWING  IIB  IIO
*
* THE FOLLOWING PARAMETERS ARE TEMPERATURE DEPENDENT AND ARE
* SIMULATED  BY THE MODEL:  ISC  VIO
*
*
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | |  | OUTPUT
*                | | |  |   | VCLAMP
*                | | |  |   |  |  GND(REFERENCE)
*                | | |  |   |  |   |
.SUBCKT HS3516   1 2 3A 4A  5     100
*
* DC PSRR FIX
Q1 11 16 13 HS3516QA
EPSRR- 16 2 TABLE {-V(4)} = (0,150U) (20,-50U)
Q2 12 15 14 HS3516QB
EPSRR+ 1 15 TABLE {V(3)} = (0,150U) (20,-50U)
*
RC1 3 11 1.447K
RC2 3 12 1.447K
C1 11 12 6.11P
RE1 13 10 1.222K
RE2 14 10 1.222K
GIEE 10 4 TABLE {V(3,4)} = (0,0) (2,0) (3,230U)
CE 10 100 0.952P
RE 10 100 869K
RP 3 4 6.289K
*
* CMRR FIX
GCM1 100 83 10 100 1
RCM1 83 84 1
LCM1 84 100 1.592U
GCM2 100 85 83 100 1
RCM2 85 86 1
LCM2 86 100 0.1592U
RCM3 86 100 10
GCM 100 21 85 100 3.087N
*
GA 21 100 11 12 691U
*
* PSRR VS FREQ FIX
GPSRR- 21 100 88 100 1
GVP- 100 88 4 100 1
RVP- 88 100 1
LVP- 88 100 0.1P
GPSRR+ 21 100 89 100 1
GVP+ 100 89 3 100 1
RVP+ 89 100 1
LVP+ 89 100 10P
*
R2 21 100 100K
C2 21 22 10P
GB 22 100 21 100 362.6
*
* VOLTAGE CLAMP
*RCL 9 100 100K
*VICL1 9 53
*VICL2 54 53
*RVOUT 54 55 10K
*EOUT 55 100 5 100 1
*WCL3 54 56 VICL3 CL
*RX 56 100 100K
*ICL+ 56 100 4M
*WCL4 54 57 VICL4 CL
*RY 57 100 100K
*ICL- 100 57 4M
*ECL1 47 100 9 100 1
*WCL1 47 48 VICL1 CL
*D8 48 49 SMX10114DD
*.MODEL SMX10114DD D (IS=1.075U)
*VICL3 49 6
*ECL2 52 100 9 100 1
*WCL2 52 51 VICL2 CL
*D9 50 51 SMX10114DE
*.MODEL SMX10114DE D (IS=15.28N)
*VICL4 6 50
*.MODEL CL ISWITCH (ION=2U IOFF=0 RON=1 ROFF=0.1MEG)
*
* END OF VCLAMP SECTION
RO2 22 100 20
D1 22 31 HS3516DA
D2 31 22 HS3516DC
EC 31 100 5 100 1.0
*
* I(VCC) FIX
RO1 22 6 30
VIOUT 6 5 0
D5 3 7 HS3516DB
R5 7 100 1MEG
F5 7 100 VIOUT 1
D6 8 4 HS3516DB
R6 8 100 1MEG
F6 8 100 VIOUT 1
*
* POWER OFF FIX
VIVP+ 3A 3
WVP+ 3 3B VIVP+ CL1
VIVP- 4 4A
WVP- 4 4B VIVP- CL1
.MODEL CL1 ISWITCH(
+        RON = 0.1
+       ROFF = 0.079MEG
+        ION = 0.5U
+       IOFF = 1N
+ )
*
* CLIPPING FIX
D3 5 24 HS3516DB
EVC 3B 24 TABLE {V(3)} = (0,0.805) (5,2.255) (10,2.305)
D4 25 5 HS3516DB
EVE 25 4B TABLE {-V(4)} = (0,0.806) (5,3.179) (10,3.226)
*
.MODEL HS3516DA D (
+         IS = 191E-12
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL HS3516DC D (
+         IS = 45.32E-12
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
F+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL HS3516DB D (
+         IS = 0.8F
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL HS3516QA NPN (
+         IS = 0.816F
+         BF = 6446
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
.MODEL HS3516QB NPN (
+         IS = 0.8F
+         BF = 9729
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
.ENDS HS3516
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LF411    1 2 3 4 5
*
  c1   11 12 4.196E-12
  c2    6  7 10.00E-12
  css  10 99 1.333E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 31.83E6 -1E3 1E3 30E6 -30E6
  ga    6  0 11 12 251.4E-6
  gcm   0  6 10 99 2.514E-9
  iss  10  4 dc 170.0E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   3 11 3.978E3
  rd2   3 12 3.978E3
  ro1   8  5 50
  ro2   7 99 25
  rp    3  4 15.00E3
  rss  10 99 1.176E6
  vb    9  0 dc 0
  vc    3 53 dc 1.500
  ve   54  4 dc 1.500
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18 Rs=1m)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=12.50E-12 Beta=743.3E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LF412    1 2 3 4 5
*
  x_lf412 1 2 3 4 5 LF411
.ends
*$
*-----------------------------------------------------------------------------
* created using Parts release 7.1p on 08/12/96 at 16:13
*
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM12     1 2 3 4 5
*
  c1   11 12 37.321E-12
  c2    6  7 20.000E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 5.0767E9 -1E3 1E3 5E9 -5E9
  ga    6  0 11 12 262.64E-6
  gcm   0  6 10 99 13.332E-9
  iee   3 10 dc 184.30E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx1
  q2   12  1 14 qx2
  r2    6  9 100.00E3
  rc1   4 11 3.8075E3
  rc2   4 12 3.8075E3
  re1  13 10 3.5207E3
  re2  14 10 3.5207E3
  ree  10 99 1.0852E6
  ro1   8  5 75.000E-3
  ro2   7 99 75.000E-3
  rp    3  4 36.004
  vb    9  0 dc 0
  vc    3 53 dc 5.6654
  ve   54  4 dc 5.6654
  vlim  7  8 dc 0
  vlp  91  0 dc 13.000E3
  vln   0 92 dc 13.000E3
.model dx D(Is=800.00E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx1 PNP(Is=800.00E-18 Bf=552.55)
.model qx2 PNP(Is=859.6504E-18 Bf=677.97)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt LM101A   1 2 3 4 5 6 7
*
  c1   11 12 8.661E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 37.73E6 -1E3 1E3 40E6 -40E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 2.988E-9
  iee  10  4 dc 15.06E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.849E3
  re2  14 10 1.849E3
  ree  10 99 13.28E6
  ro1   8  5 50
  ro2   7 99 25
  rp    3  4 15.11E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=250)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt LM108    1 2 3 4 5 6 7
*
  c1   11 12 5.460E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 83.87E6 -1E3 1E3 80E6 -80E6
  ga    6  0 11 12 150.8E-6
  gcm   0  6 10 99 1.508E-9
  iee  10  4 dc 18.00E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 6.631E3
  rc2   3 12 6.631E3
  re1  13 10 3.757E3
  re2  14 10 3.757E3
  ree  10 99 11.11E6
  ro1   8  5 50
  ro2   7 99 25
  rp    3  4 106.4E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 6
  vln   0 92 dc 6
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=11.25E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM118    1 2 3 4 5
*
  c1   11 12 2.887E-12
  c2    6  7 20.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 636.5E3 -1E3 1E3 600E3 -600E3
  ga    6  0 11 12 12.57E-3
  gcm   0  6 10 99 125.7E-9
  iee  10  4 dc 1.400E-3
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 79.57
  rc2   3 12 79.57
  re1  13 10 42.61
  re2  14 10 42.61
  ree  10 99 142.8E3
  ro1   8  5 50
  ro2   7 99 25
  rp    3  4 9.678E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 22
  vln   0 92 dc 22
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=5.833E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM124    1 2 3 4 5
*
  c1   11 12 2.887E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 21.22E6 -1E3 1E3 20E6 -20E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 10.60E-9
  iee   3 10 dc 15.09E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   4 11 5.305E3
  rc2   4 12 5.305E3
  re1  13 10 1.845E3
  re2  14 10 1.845E3
  ree  10 99 13.25E6
  ro1   8  5 50
  ro2   7 99 25
  rp    3  4 9.082E3
  vb    9  0 dc 0
  vc    3 53 dc 1.500
  ve   54  4 dc 0.65
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx PNP(Is=800.0E-18 Bf=166.7)
.ends
*$
*
* MANUFACTURERS PART NO. = LM124W  (TEXAS INSTRUMENTS)
* SUBTYPE: OP_AMP
* THIS FILE CONTAINS A PRE-RAD MODEL OF THE LM124
* WHICH HAS BEEN VERIFIED FOR USE WITH A .TEMP CARD.
* THIS MODEL MAY BE USED FOR ALL OF THE FOLLOWING DEVICES :
* LM124
* LM124J
* LM124W
*
* THE FOLLOWING MODEL WAS DERIVED USING MEASURED DATA.
*
* THIS MODEL CAN BE USED WITH A .TEMP CARD OVER THE TEMPERATURE RANGE
* OF -55 C TO 125 C.
* THE FOLLOWING PARAMETERS ARE INSENSITIVE TO TEMPERATURE CHANGES AND
* ARE  SIMULATED ACCURATELY BY THE MODEL: CMRR  GAIN  PSRR  OUTPUT
* VOLTAGE SWING  HIGH LEVEL ONLY
*
* THE FOLLOWING PARAMETERS ARE NOT SIMULATED BY THE MODEL OVER
* TEMPERATURE:  IIB   ICC   GBW   OUTPUT VOLTAGE SWING LOW LEVEL
*
* THIS MODEL DOES NOT SIMULATE VOS (INPUT OFFSET VOLTAGE) OR IOS (INPUT
* OFFSET  CURRENT).
*
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | | GND(REFERENCE)
.SUBCKT LM124A   1 2 3 4 5  100
*
C1   11 12 2.887E-12
C2    6  7 30.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  100 POLY(2) (3,100) (4,100) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 21.22E6 -20E6 20E6 20E6 -20E6
GA    6  100 11 12 188.5E-6
GCM   100  6 10 99 10.60E-9
IEE   3 10 DC 15.09E-6
HLIM 90  100 VLIM 1K
Q1   11  2 13 QX
Q2   12  1 14 QX
R2    6  9 100.0E3
RC1   4 11 5.305E3
RC2   4 12 5.305E3
RE1  13 10 1.845E3
RE2  14 10 1.845E3
REE  10 99 13.25E6
RO1   8  5 50
RO2   7 99 25
RP    3  4 9.082E3
VB    9  100 DC 0
VC    3 53 DC 1.500
VE   54  4 DC 0
VLIM  7  8 DC 0
VLP  91  100 DC 40
VLN   100 92 DC 40
.MODEL DX D(
+         IS = 800.0E-18
+         RS = 1
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.MODEL QX PNP(
+         IS = 800.0E-18
+         BF = 166.7
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.ENDS
*$
*
* MANUFACTURERS PART NO. = LM124W  (TEXAS INSTRUMENTS)
* SUBTYPE: OP_AMP
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT MODEL OF THE LM124.
* THIS MODEL MAY BE USED FOR ALL OF THE FOLLOWING DEVICES :
* LM124
* LM124J
* LM124W
*
*
* IT MODELS POWER-UP, POWER-DOWN, AND POWER OFF CONDITIONS,
* SINGLE SUPPLY APPLICATIONS, AC PSRR, DC PSRR, AC CMRR, VSAT, IIB, IIO,
* VIO, ISC, SR, PM, GBP, ICC, AND RO(AC).
*-----------------------------------------------------------------------------
*-----------------------------------------------------------------------------
* THE FOLLOWING SPECIFICATIONS ARE SIMULATED IN THE MODEL FOR +/-15 V
* SUPPLIES:
*  VIO = -2.05 MV, VSAT = +13.6 V, VSAT- = -14.3 V, IB = 15.2 NA, IIO = 1 NA
*  GBP = 0.91M HZ, PM = 49 DEG, CMRR = 87 DB, RO(AC) = 31 OHMS, ISC+ = 40 MA
*  ISC- = -20 MA, SR+ = 0.3 V/US, SR- = -0.33 V/US
*
* MODIFIED SPECS:
* DC PSRR = 108 DB, AC PSRR MODELED; ISUPPLY = IBIAS + ILOAD, VSAT VARIES WITH
* SUPPLY VOLTAGES, ALSO MODELS SINGLE SUPPLY APPLICATIONS; E.G. VCC+ = 5 V,
* VCC- = 0 V, VSAT+ = 3 V, VSAT- = 5 MV; POWER NOT CONNECTED MODELED; POWER-
* UP AND POWER-DOWN MODELED.
*
* THIS MODEL CAN BE USED WITH A .TEMP CARD OVER THE TEMPERATURE RANGE
* OF  -55 C TO 125 C.
*
* THE FOLLOWING PARAMETERS ARE INSENSITIVE TO TEMPERATURE CHANGES AND
* ARE SIMULATED ACCURATELY BY THE MODEL: CMRR  GAIN  ICC  PSRR  SR
* OVERDRIVE  RECOVERY TIME   OUTPUT VOLTAGE SWING  IIB  IIO
*
* THE FOLLOWING PARAMETERS ARE TEMPERATURE DEPENDENT AND ARE
* SIMULATED  BY THE MODEL:  ISC  VIO
*
*
* CONNECTIONS:        NON-INVERTING INPUT
*                     | INVERTING INPUT
*                     | | POSITIVE POWER SUPPLY
*                     | | | NEGATIVE POWER SUPPLY
*                     | | |  | OUTPUT
*                     | | |  |  |  GND(REFERENCE)
.SUBCKT LM124/TEMP    1 2 3A 4A 5  100
*
* DC PSRR FIX
Q1 11 16 13 LM124QA
EPSRR- 16 2 TABLE {-V(4)} = (0,622U) (16,-41.45U)
Q2 12 15 14 LM124QB
EPSRR+ 1 15 TABLE {V(3)} = (0,552U) (16,-36.82U)
*
RC1 4 11 16.182K
RC2 4 12 16.182K
C1 11 12 5.71P
RE1 13 10 467
RE2 14 10 467
GIEE 3 10 TABLE {V(3,4)} = (0,0) (2,0) (3 3.291U)
CE 10 100 0.661P
RE 10 100 60.77MEG
*
* SUPPLY CURRENT FOR 1/4 CURRENT OF IC.
* PLACE AN RP IN PARALLEL FOR EACH UNUSED OPAMP ON IC.
RP 3 4 80.7K
*
* CMRR FIX
GCM1 100 83 10 100 1
RCM1 83 84 1
LCM1 84 100 15.92U
GCM2 100 85 83 100 1
RCM2 85 86 1
LCM2 86 100 1.592U
RCM3 86 100 10
GCM 100 21 85 100 2.63N
*
GA 21 100 11 12 61.797U
*
* PSRR VS FREQ FIX
GPSRR- 21 100 88 100 1
GVP- 100 88 4 100 1
RVP- 88 100 1
LVP- 88 100 10P
GPSRR+ 21 100 89 100 1
GVP+ 100 89 3 100 1
RVP+ 89 100 1
LVP+ 89 100 0.1P
*
R2 21 100 100K
C2 21 22 10P
GB 22 100 21 100 777.93
RO2 22 100 80
D1 22 31 LM124DA
D2 31 22 LM124DC
EC 31 100 5 100 1.0
*
* I(VCC) FIX
RO1 22 6 31
VIOUT 6 5 0
D5 3 7 LM124DB
R5 7 100 1MEG
F5 7 100 VIOUT 1
D6 8 4 LM124DB
R6 8 100 1MEG
F6 8 100 VIOUT 1
*
* POWER OFF FIX
VIVP+ 3A 3
WVP+ 3 3B VIVP+ CL1
VIVP- 4 4A
WVP- 4 4B VIVP- CL1
.MODEL CL1 ISWITCH(
+        RON = 0.1
+       ROFF = 18MEG
+        ION = 0.5U
+       IOFF = 1N
+ )
*
* CLIPPING FIX
D3 5 24 LM124DB
EVC 3B 24 TABLE {V(3)} = (0,0.815) (5,2.115) (10,2.115) (16,2.235)
D4 25 5 LM124DB
EVE 25 4B TABLE {-V(4)} = (0,0.798) (5,1.498) (16,1.498)
*
.MODEL LM124DA D (
+         IS = 383E-21
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL LM124DC D (
+         IS = 9.907N
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL LM124DB D (
+         IS = 0.8F
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL LM124QA PNP (
+         IS = 0.8666F
+         BF = 111.7
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
.MODEL LM124QB PNP (
+         IS = 0.8F
+         BF = 104.6
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
.ENDS
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM158    1 2 3 4 5
*
  x_lm158 1 2 3 4 5 LM124
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt LM201A   1 2 3 4 5 6 7
*
  x_lm201a 1 2 3 4 5 6 7 LM101A
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt LM208    1 2 3 4 5 6 7
*
  x_lm208 1 2 3 4 5 6 7 LM108
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM218    1 2 3 4 5
*
  x_lm218 1 2 3 4 5 LM118
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM224    1 2 3 4 5
*
  x_lm224 1 2 3 4 5 LM124
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM258    1 2 3 4 5
*
  x_lm258 1 2 3 4 5 LM124
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt LM301A   1 2 3 4 5 6 7
*
  c1   11 12 8.661E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 21.22E6 -1E3 1E3 20E6 -20E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.14E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.839E3
  re2  14 10 1.839E3
  ree  10 99 13.21E6
  ro1   8  5 50
  ro2   7 99 25
  rp    3  4 15.11E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=107.1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt LM308    1 2 3 4 5 6 7
*
  c1   11 12 5.460E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 83.87E6 -1E3 1E3 80E6 -80E6
  ga    6  0 11 12 150.8E-6
  gcm   0  6 10 99 1.508E-9
  iee  10  4 dc 18.00E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 6.631E3
  rc2   3 12 6.631E3
  re1  13 10 3.756E3
  re2  14 10 3.756E3
  ree  10 99 11.11E6
  ro1   8  5 50
  ro2   7 99 25
  rp    3  4 106.4E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 6
  vln   0 92 dc 6
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=6.000E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM318    1 2 3 4 5
*
  c1   11 12 2.887E-12
  c2    6  7 20.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 636.5E3 -1E3 1E3 600E3 -600E3
  ga    6  0 11 12 12.57E-3
  gcm   0  6 10 99 125.7E-9
  iee  10  4 dc 1.400E-3
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 79.57
  rc2   3 12 79.57
  re1  13 10 42.61
  re2  14 10 42.61
  ree  10 99 142.8E3
  ro1   8  5 50
  ro2   7 99 25
  rp    3  4 9.678E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 22
  vln   0 92 dc 22
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=4.667E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM324    1 2 3 4 5
*
  c1   11 12 2.887E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 21.22E6 -1E3 1E3 20E6 -20E6

  fpos a 0 vlim 1
  w2 3 a vlim sw2
  .model sw2 iswitch (ron=1 ion=0 ioff=-1u roff=10meg)
  w1 a 0 vlim sw1
  .model sw1 iswitch (roff=10meg ioff=0 ion=-1u ron=1)

  fneg 0 b vlim -1
  w3 4 b vlim sw3
  .model sw3 iswitch (ron=1 ion=-1u ioff=0 roff=10meg)
  w4 b 0 vlim sw4
  .model sw4 iswitch (roff=10meg ioff=-1u ion=0 ron=1)


  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 59.61E-9
  iee   3 10 dc 15.09E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   4 11 5.305E3
  rc2   4 12 5.305E3
  re1  13 10 1.845E3
  re2  14 10 1.845E3
  ree  10 99 13.25E6
  ro1   8  5 50
  ro2   7 99 25
  rp    3  4 9.082E3
  vb    9  0 dc 0
  vc    3 53 dc 1.500
  ve   54  4 dc 0.65
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx PNP(Is=800.0E-18 Bf=166.7)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM358    1 2 3 4 5
*
  x_lm358 1 2 3 4 5 LM324
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt lm675    1 2 3 4 5
*
  c1   11 12 8.660E-12
  c2    6  7 15.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 7.717E9 -1E3 1E3 7E9 -7E9
  ga    6  0 11 12 518.4E-6
  gcm   0  6 10 99 16.40E-9
  iee   3 10 dc 120.4E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   4 11 1.929E3
  rc2   4 12 1.929E3
  re1  13 10 1.493E3
  re2  14 10 1.493E3
  ree  10 99 1.661E6
  ro1   8  5 50.00E-3
  ro2   7 99 50.00E-3
  rp    3  4 2.796E3
  vb    9  0 dc 0
  vc    3 53 dc 4
  ve   54  4 dc 4
  vlim  7  8 dc 0
  vlp  91  0 dc 3.000E3
  vln   0 92 dc 3.000E3
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx PNP(Is=800.0E-18 Bf=300)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt LM709    1 2 3 4 5 6 7
  x_lm709 1 2 3 4 5 6 7 uA709
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt lm709a   1 2 3 4 5 6 7
*
  c1   11 12 8.660E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 716.2E3 -1E3 1E3 720E3 -720E3
  ga    6  0 11 12 1.257E-3
  gcm   0  6 10 99 3.974E-9
  iee  10  4 dc 100.2E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 795.8
  rc2   3 12 795.8
  re1  13 10 277.9
  re2  14 10 277.9
  ree  10 99 1.996E6
  ro1   8  5 50
  ro2   7 99 50
  rp    3  4 12.50E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 42
  vln   0 92 dc 42
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=500)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt lm709c   1 2 3 4 5 6 7
*
  c1   11 12 8.660E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 716.2E3 -1E3 1E3 720E3 -720E3
  ga    6  0 11 12 1.257E-3
  gcm   0  6 10 99 39.74E-9
  iee  10  4 dc 100.6E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 795.8
  rc2   3 12 795.8
  re1  13 10 276.8
  re2  14 10 276.8
  ree  10 99 1.988E6
  ro1   8  5 50
  ro2   7 99 50
  rp    3  4 11.69E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 42
  vln   0 92 dc 42
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=166.7)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM741    1 2 3 4 5
*
  x_lm741 1 2 3 4 5 uA741
.ends
*$
*----------------------------------------------------------------------------
* created using Parts release 7.1p on 07/24/96 at 15:00
*
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt LM759C   1 2 3 4 5
*
  c1   11 12 5.6383E-12
  c2    6  7 12.000E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 76.126E6 -1E3 1E3 76E6 -76E6
  ga    6  0 11 12 101.41E-6
  gcm   0  6 10 99 1.0187E-9
  iee   3 10 dc 6.4604E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx1
  q2   12  1 14 qx2
  r2    6  9 100.00E3
  rc1   4 11 9.8609E3
  rc2   4 12 9.8609E3
  re1  13 10 1.7008E3
  re2  14 10 1.7008E3
  ree  10 99 30.958E6
  ro1   8  5 5
  ro2   7 99 5
  rp    3  4 2.5013E3
  vb    9  0 dc 0
  vc    3 53 dc 3.0212
  ve   54  4 dc 3.0212
  vlim  7  8 dc 0
  vlp  91  0 dc 500
  vln   0 92 dc 500
.model dx D(Is=800.00E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx1 PNP(Is=800.00E-18 Bf=59.618)
.model qx2 PNP(Is=831.5365E-18 Bf=67.616)
.ends
*$
*-----------------------------------------------------------------------------
* created using Parts release 7.1p on 07/25/96 at 15:01
*
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt MAX402   1 2 3 4 5
*
  c1   11 12 10.118E-12
  c2    6  7 30.000E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 58.987E3 -1E3 1E3 59E3 -59E3
  ga    6  0 11 12 446.73E-6
  gcm   0  6 10 99 7.9511E-9
  iee   3 10 dc 219.00E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx1
  q2   12  1 14 qx2
  r2    6  9 100.00E3
  rc1   4 11 2.2385E3
  rc2   4 12 2.2385E3
  re1  13 10 2.0022E3
  re2  14 10 2.0022E3
  ree  10 99 913.23E3
  ro1   8  5 222
  ro2   7 99 222
  rp    3  4 268.23
  vb    9  0 dc 0
  vc    3 53 dc 1.7178
  ve   54  4 dc 1.7178
  vlim  7  8 dc 0
  vlp  91  0 dc 3.5000
  vln   0 92 dc 3.5000
.model dx D(Is=800.00E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx1 PNP(Is=800.00E-18 Bf=51.859E3)
.model qx2 PNP(Is=815.6159E-18 Bf=57.375E3)
.ends
*$
*-----------------------------------------------------------------------------
* created using Parts release 7.1p on 08/12/96 at 09:51
*
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt MAX403   1 2 3 4 5
*
  c1   11 12 10.503E-12
  c2    6  7 30.000E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 117.50E3 -1E3 1E3 120E3 -120E3
  ga    6  0 11 12 2.2619E-3
  gcm   0  6 10 99 226.19E-9
  iee   3 10 dc 1.2510E-3
  hlim 90  0 vlim 1K
  q1   11  2 13 qx1
  q2   12  1 14 qx2
  r2    6  9 100.00E3
  rc1   4 11 442.10
  rc2   4 12 442.10
  re1  13 10 400.74
  re2  14 10 400.74
  ree  10 99 159.87E3
  ro1   8  5 38
  ro2   7 99 38
  rp    3  4 275.87
  vb    9  0 dc 0
  vc    3 53 dc 1.7941
  ve   54  4 dc 1.7941
  vlim  7  8 dc 0
  vlp  91  0 dc 2.5000
  vln   0 92 dc 2.5000
.model dx D(Is=800.00E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx1 PNP(Is=800.00E-18 Bf=59.261E3)
.model qx2 PNP(Is=812.4685E-18 Bf=65.532E3)
.ends
*$
*-----------------------------------------------------------------------------
* created using Parts release 7.1p on 08/29/96 at 16:15
*
* connections:     input
*                  |  adjustment pin
*                  |  |   output
*                  |  |   |
.SUBCKT LM317     IN ADJ OUT
*
* POSITIVE ADJUSTABLE VOLTAGE REGULATOR
*
JADJ IN ADJ ADJ JADJMOD ;ADJUSTMENT PIN CURRENT
VREF 4 ADJ 1.250
DBK IN 13 DMOD
*
* ZERO OF RIPPLE REJECTION
*
*
*
CBC 13 15 800.0E-12
RBC 15 5 1.000E3
*
QPASS 13 5 OUT QPASSMOD
RB1 7 6 1
RB2 6 5 128.3
*
* CURRENT LIMITING
*
DSC 6 11 DMOD
ESC 11 OUT VALUE={5.646-.6667*V(6,5)*V(13,5)}
*
* FOLDBACK CURRENT
*
DFB 6 12 DMOD
EFB 12 OUT VALUE={8.822-.4024*V(13,5)+5.250E-3*V(13,5)*V(13,5)
+ -.6667*V(13,5)*V(6,5)}
*
EB 7 OUT 8 OUT 6.939
*
* ZERO OF OUTPUT IMPEDANCE
*
RP 9 8 100
CPZ 10 OUT 3.183E-6
*
DPU 10 OUT DMOD ;POWER-UP CLAMPLING DIODE
RZ 8 10 .1
EP 9 OUT 4 OUT 100
RI OUT 4 100MEG
*
.MODEL QPASSMOD NPN (IS=30F BF=50 VAF=1.500 NF=1.701)
.MODEL JADJMOD NJF (BETA=50.00E-6 VTO=-1)
.MODEL DMOD D (IS=30F N=1.701)
.ENDS
*$
*-----------------------------------------------------------------------------
* created using Parts release 7.1p on 08/26/96 at 10:12
*
* connections:    Anode
*                 |  Cathode
*                 |  |
.SUBCKT LM385     A  K
*
* TWO-TERMINAL VOLTAGE REFERENCE
*
DFWD A K DF
GREV A K VALUE={LIMIT(20.00E-3*(EXP(V(A,K)/5.682E3)-1),-10M,0)}
RZ A 1 .102
GZ 2 1 VALUE={LIMIT(EXP(V(2,1)/198.0E-6),0,20.00E-3)}
EBV K 2 3 0 1
RBV 3 0 1.237E3 TC=1.139E-6 -346.8E-9
IBV 0 3 DC 1M
*
.MODEL DF D(IS=39.12E-15 RS=12.18 IKF=0 N=.9983 XTI=3)
.ENDS
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt mc1458   1 2 3 4 5
*
  c1   11 12 8.660E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 42.44E6 -1E3 1E3 42E6 -42E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.837E3
  re2  14 10 1.837E3
  ree  10 99 13.19E6
  ro1   8  5 25
  ro2   7 99 25
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 20
  vln   0 92 dc 20
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt mc1458c  1 2 3 4 5
*
  c1   11 12 8.660E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 42.44E6 -1E3 1E3 42E6 -42E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.837E3
  re2  14 10 1.837E3
  ree  10 99 13.19E6
  ro1   8  5 25
  ro2   7 99 25
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 20
  vln   0 92 dc 20
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt mc1458s  1 2 3 4 5
*
  c1   11 12 8.660E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 42.44E6 -1E3 1E3 42E6 -42E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 600.4E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 5.215E3
  re2  14 10 5.215E3
  ree  10 99 333.1E3
  ro1   8  5 25
  ro2   7 99 25
  rp    3  4 28.13E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 20
  vln   0 92 dc 20
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=1.500E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt mc1558   1 2 3 4 5
*
  c1   11 12 8.660E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 42.44E6 -1E3 1E3 42E6 -42E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.837E3
  re2  14 10 1.837E3
  ree  10 99 13.19E6
  ro1   8  5 25
  ro2   7 99 25
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 20
  vln   0 92 dc 20
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt mc1558s  1 2 3 4 5
*
  c1   11 12 8.660E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 42.44E6 -1E3 1E3 42E6 -42E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 600.4E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 5.215E3
  re2  14 10 5.215E3
  ree  10 99 333.1E3
  ro1   8  5 25
  ro2   7 99 25
  rp    3  4 28.13E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 20
  vln   0 92 dc 20
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=1.500E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt mc1709   1 2 3 4 5 6 7
*
  c1   11 12 8.660E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 716.2E3 -1E3 1E3 720E3 -720E3
  ga    6  0 11 12 1.257E-3
  gcm   0  6 10 99 39.74E-9
  iee  10  4 dc 100.4E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 795.8
  rc2   3 12 795.8
  re1  13 10 277.4
  re2  14 10 277.4
  ree  10 99 1.992E6
  ro1   8  5 50
  ro2   7 99 50
  rp    3  4 11.69E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=250)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt mc1709a  1 2 3 4 5 6 7
*
  c1   11 12 8.660E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 716.2E3 -1E3 1E3 720E3 -720E3
  ga    6  0 11 12 1.257E-3
  gcm   0  6 10 99 3.974E-9
  iee  10  4 dc 100.2E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 795.8
  rc2   3 12 795.8
  re1  13 10 277.9
  re2  14 10 277.9
  ree  10 99 1.996E6
  ro1   8  5 50
  ro2   7 99 50
  rp    3  4 12.50E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=500)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt mc1709c  1 2 3 4 5 6 7
*
  c1   11 12 8.660E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 716.2E3 -1E3 1E3 720E3 -720E3
  ga    6  0 11 12 1.257E-3
  gcm   0  6 10 99 39.74E-9
  iee  10  4 dc 100.6E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 795.8
  rc2   3 12 795.8
  re1  13 10 276.8
  re2  14 10 276.8
  ree  10 99 1.988E6
  ro1   8  5 50
  ro2   7 99 50
  rp    3  4 11.69E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=166.7)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt mc1741   1 2 3 4 5
*
  c1   11 12 8.660E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 42.44E6 -1E3 1E3 42E6 -42E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.837E3
  re2  14 10 1.837E3
  ree  10 99 13.19E6
  ro1   8  5 25
  ro2   7 99 25
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 20
  vln   0 92 dc 20
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt mc33076  1 2 3 4 5
*
  c1   11 12 11.72E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 6.063E6 -1E3 1E3 6E6 -6E6
  ga    6  0 11 12 659.7E-6
  gcm   0  6 10 99 20.86E-9
  iee   3 10 dc 78.20E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   4 11 1.516E3
  rc2   4 12 1.516E3
  re1  13 10 850.4
  re2  14 10 850.4
  ree  10 99 2.558E6
  ro1   8  5 50
  ro2   7 99 50
  rp    3  4 10.89E3
  vb    9  0 dc 0
  vc    3 53 dc 1.200
  ve   54  4 dc 1.200
  vlim  7  8 dc 0
  vlp  91  0 dc 250
  vln   0 92 dc 250
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx PNP(Is=800.0E-18 Bf=390)
.ends
*$
*
* MANUFACTURERS PART NO. = SMX10114
* SUBTYPE: OP_AMP
* THIS FILE CONTAINS A PRE-RAD MODEL.  IT HAS BEEN VERIFIED FOR USE WITH A
* .TEMP CARD.  COMMENTS CONCERNING VALIDITY ARE IN THE SECTION PRECEEDING
* THE MODEL.
*
* THIS MODEL CAN BE USED WITH A .TEMP CARD OVER THE TEMPERATURE RANGE
* OF  -55 C TO 125 C.
*
* THE FOLLOWING PARAMETERS ARE INSENSITIVE TO TEMPERATURE CHANGES AND
* ARE  SIMULATED ACCURATELY BY THE MODEL: CMRR  GAIN  PSRR  OUTPUT
* VOLTAGE SWING
*
* THE FOLLOWING PARAMETERS ARE TEMPERATURE DEPENDENT BUT ARE NOT
* SIMULATED  BY THE MODEL: IIB  ISC  TOR  SR  ICC
*
* ALL ARE WITHIN THE PRODUCT SPEC LIMITS OVER TEMPERATURE.
*
* THIS MODEL DOES NOT SIMULATE VOS (INPUT OFFSET VOLTAGE) OR IOS (INPUT
* OFFSET  CURRENT).  IT DOES CORRECTLY SIMULATE PHASE MARGIN, UNITY GAIN
* BANDWIDTH,  CMRR, MAX. POSITIVE AND NEGATIVE OUTPUT VOLTAGE SWING (ONLY
* WITH SYMMETRIC POWER SUPPLIES),  POWER DISSIPATION, AND FREQUENCY
* RESPONSE(PHASE LAG ABOVE  100HZ & GAIN ABOVE 10HZ).
*
*
*
*
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |  GND(REFERENCE)
.SUBCKT MPR155   1 2 3 4 5  100
*
C1   11 12 4.502E-12
C2    6  7 10.00E-12
CSS  10 99 2.727E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  100 POLY(2) (3,100) (4,100) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 2.809E6 -3E6 3E6 3E6 -3E6
GA    6  100 11 12 565.5E-6
GCM   100  6 10 99 5.655E-9
ISS   3 10 DC 280.0E-6
HLIM 90  100 VLIM 1K
J1   11  2 10 JX
J2   12  1 10 JX
R2    6  9 100.0E3
RD1   4 11 1.768E3
RD2   4 12 1.768E3
RO1   8  5 50
RO2   7 99 25
RP    3  4 7.500E3
RSS  10 99 714.3E3
VB    9  100 DC 0
VC    3 53 DC 2
VE   54  4 DC 2.500
VLIM  7  8 DC 0
VLP  91  100 DC 45
VLN   100 92 DC 45
.MODEL DX D(
+         IS = 800.0E-18
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+ )
.MODEL JX PJF(
+        VTO = -1
+       BETA = 2.284E-3
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CGS = 0
+        CGD = 0
+         PB = 1
+         IS = 5.000E-12
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.ENDS MPR155
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt OP-07    1 2 3 4 5
*
  c1   11 12 8.661E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 221.0E6 -1E3 1E3 200E6 -200E6
  ga    6  0 11 12 113.1E-6
  gcm   0  6 10 99 56.69E-12
  iee  10  4 dc 6.002E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 8.841E3
  rc2   3 12 8.841E3
  re1  13 10 219.4
  re2  14 10 219.4
  ree  10 99 33.32E6
  ro1   8  5 40
  ro2   7 99 20
  rp    3  4 12.03E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 30
  vln   0 92 dc 30
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=3.000E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt OP-27    1 2 3 4 5
*
  c1   11 12 5.460E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 39.78E6 -1E3 1E3 40E6 -40E6
  ga    6  0 11 12 1.508E-3
  gcm   0  6 10 99 755.9E-12
  iee  10  4 dc 84.02E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 663.1
  rc2   3 12 663.1
  re1  13 10 47.24
  re2  14 10 47.24
  ree  10 99 2.380E6
  ro1   8  5 40
  ro2   7 99 30
  rp    3  4 9.233E3
  vb    9  0 dc 0
  vc    3 53 dc 1.200
  ve   54  4 dc 1.200
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=4.200E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt op-471a  1 2 3 4 5
*
  c1   11 12 9.741E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 9.174E9 -1E3 1E3 9E9 -9E9
  ga    6  0 11 12 1.225E-3
  gcm   0  6 10 99 1.225E-9
  iee  10  4 dc 240.0E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 816.2
  rc2   3 12 816.2
  re1  13 10 600.6
  re2  14 10 600.6
  ree  10 99 833.2E3
  ro1   8  5 50.00E-3
  ro2   7 99 50.00E-3
  rp    3  4 14.56E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=7.500E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt op-471e  1 2 3 4 5
*
  c1   11 12 9.741E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 9.174E9 -1E3 1E3 9E9 -9E9
  ga    6  0 11 12 1.225E-3
  gcm   0  6 10 99 2.180E-9
  iee  10  4 dc 240.0E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 816.2
  rc2   3 12 816.2
  re1  13 10 600.6
  re2  14 10 600.6
  ree  10 99 833.2E3
  ro1   8  5 50.00E-3
  ro2   7 99 50.00E-3
  rp    3  4 14.56E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=9.231E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt OP-471F  1 2 3 4 5
*
  c1   11 12 9.741E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 9.174E9 -1E3 1E3 9E9 -9E9
  ga    6  0 11 12 1.225E-3
  gcm   0  6 10 99 3.877E-9
  iee  10  4 dc 240.0E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 816.2
  rc2   3 12 816.2
  re1  13 10 600.6
  re2  14 10 600.6
  ree  10 99 833.2E3
  ro1   8  5 50.00E-3
  ro2   7 99 50.00E-3
  rp    3  4 14.56E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=8.000E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt OP-471G  1 2 3 4 5
*
  c1   11 12 9.741E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 9.174E9 -1E3 1E3 9E9 -9E9
  ga    6  0 11 12 1.225E-3
  gcm   0  6 10 99 3.877E-9
  iee  10  4 dc 240.1E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 816.2
  rc2   3 12 816.2
  re1  13 10 600.4
  re2  14 10 600.4
  ree  10 99 833.1E3
  ro1   8  5 50.00E-3
  ro2   7 99 50.00E-3
  rp    3  4 14.56E3
  vb    9  0 dc 0
  vc    3 53 dc 2
  ve   54  4 dc 2
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=3.000E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt OPA3581J 1 2 3 4 5
*
  c1   11 12 2.887E-12
  c2    6  7 10.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 5.029E9 -1E3 1E3 5E9 -5E9
  ga    6  0 11 12 251.3E-6
  gcm   0  6 10 99 795.3E-12
  iss  10  4 dc 200.0E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   3 11 3.979E3
  rd2   3 12 3.979E3
  ro1   8  5 .25
  ro2   7 99 .25
  rp    3  4 16.00E3
  rss  10 99 1.000E6
  vb    9  0 dc 0
  vc    3 53 dc 5
  ve   54  4 dc 5
  vlim  7  8 dc 0
  vlp  91  0 dc 50
  vln   0 92 dc 50
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=10.00E-12 Beta=315.8E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt OPA3582J 1 2 3 4 5
*
  c1   11 12 2.887E-12
  c2    6  7 10.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 15.92E9 -1E3 1E3 16E9 -16E9
  ga    6  0 11 12 251.3E-6
  gcm   0  6 10 99 795.3E-12
  iss  10  4 dc 200.0E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   3 11 3.979E3
  rd2   3 12 3.979E3
  ro1   8  5 .25
  ro2   7 99 .25
  rp    3  4 21.54E3
  rss  10 99 1.000E6
  vb    9  0 dc 0
  vc    3 53 dc 5
  ve   54  4 dc 5
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=10.00E-12 Beta=315.8E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt opa3583  1 2 3 4 5
*
  c1   11 12 2.887E-12
  c2    6  7 10.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 12.73E9 -1E3 1E3 13E9 -13E9
  ga    6  0 11 12 251.3E-6
  gcm   0  6 10 99 795.3E-12
  iss  10  4 dc 300.0E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   3 11 3.979E3
  rd2   3 12 3.979E3
  ro1   8  5 .25
  ro2   7 99 .25
  rp    3  4 35.29E3
  rss  10 99 666.7E3
  vb    9  0 dc 0
  vc    3 53 dc 10
  ve   54  4 dc 10
  vlim  7  8 dc 0
  vlp  91  0 dc 100
  vln   0 92 dc 100
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=10.00E-12 Beta=210.6E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt OPA3584J 1 2 3 4 5
*
  c1   11 12 8.727E-15
  c2    6  7 10.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 169.8E9 -1E3 1E3 170E9 -170E9
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 596.5E-12
  iss  10  4 dc 1.500E-3
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   3 11 5.305E3
  rd2   3 12 5.305E3
  ro1   8  5 .25
  ro2   7 99 .25
  rp    3  4 46.15E3
  rss  10 99 133.3E3
  vb    9  0 dc 0
  vc    3 53 dc 5
  ve   54  4 dc 5
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=10.00E-12 Beta=23.69E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:    non-inverting input
*                 | inverting input
*                 | | positive power supply
*                 | | | negative power supply
*                 | | | | output
*                 | | | | |
.subckt pm-741    1 2 3 4 5
*
  c1   11 12 8.660E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 42.44E6 -1E3 1E3 42E6 -42E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.837E3
  re2  14 10 1.837E3
  ree  10 99 13.19E6
  ro1   8  5 25
  ro2   7 99 25
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 20
  vln   0 92 dc 20
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
*$
*
* MANUFACTURERS PART NO. = SMX10114  (TEXAS INSTRUMENTS)
* SUBTYPE: OP_AMP
* THIS FILE CONTAINS A PRE-RAD MODEL WHICH HAS BEEN VERIFIED
* FOR USE WITH A .TEMP CARD.  COMMENTS CONCERNING VALIDITY ARE IN THE
* SECTION  PRECEDING THE MODEL.
*
* IT MODELS POWER-UP, POWER-DOWN, AND POWER OFF CONDITIONS,
* SINGLE SUPPLY APPLICATIONS, AC PSRR, DC PSRR, AC CMRR, VSAT, IIB, IIO,
* VIO, ISC, SR, PM, GBP, ICC, AND RO(AC). THE VOLTAGE CLAMPING PIN HAS
* BEEN MODELED. IT HAS BEEN COMMENTED OUT WITH THE * SYMBOL BECAUSE IT
* CAN  CAUSE CONVERGENCE PROBLEMS. TO ADD TO THE MODEL ADD PIN 9 ON THE
* .SUBCKT  LINE AND REMOVE THE * FROM THE LINES DEFINING THE CLAMP PIN IN
* THE MODEL.  IF IT CAUSES A CONVERGENCE PROBLEM USE ITL4=300 IN THE
* .OPTION STATEMENT.

*
*
*-----------------------------------------------------------------------------
* THE FOLLOWING SPECIFICATIONS ARE SIMULATED IN THE MODEL FOR +/-15 V
* SUPPLIES:
*  VIO = 1.13 MV, VSAT = +13.54 V, VSAT- = -13.5 V, IB = 94.5 PA, IIO = 49 PA
*  GBP = 9.5MHZ, PM = 55.3 DEG, CMRR = 81.2 DB, RO(AC) = 19 OHMS, ISC+ = 44 MA
*  ISC- = -28 MA, SR+ = 22 V/US, SR- = -61.5 V/US
*
* MODIFIED SPECS:
* DC PSRR = 100 DB, AC PSRR MODELED; ISUPPLY = IBIAS + ILOAD, VSAT VARIES WITH
* SUPPLY VOLTAGES, ALSO MODELS SINGLE SUPPLY APPLICATIONS; E.G. VCC+ = 5 V,
* VCC- = 0 V, VSAT+ = 3 V, VSAT- = 5 MV; POWER NOT CONNECTED MODELED; POWER-
* UP  AND POWER-DOWN MODELED. ERRORS IN IB AND IIO DUE TO GMIN ARE FIXED.
*
* THIS MODEL CAN BE USED WITH A .TEMP CARD OVER THE TEMPERATURE RANGE
* OF  -55 C TO 125 C.
*
* THE FOLLOWING PARAMETERS ARE INSENSITIVE TO TEMPERATURE CHANGES AND
* ARE  SIMULATED ACCURATELY BY THE MODEL: CMRR  GAIN  ICC  PSRR  SR
* OVERDRIVE RECOVERY TIME   OUTPUT VOLTAGE SWING  IIB  IIO
*
* THE FOLLOWING PARAMETERS ARE TEMPERATURE DEPENDENT AND ARE
* SIMULATED  BY THE MODEL:  ISC  VIO
*
*
* CONNECTIONS:   NON-INVERTING INPUT
*                 | INVERTING INPUT
*                 | | POSITIVE POWER SUPPLY
*                 | | | NEGATIVE POWER SUPPLY
*                 | | |  | OUTPUT
*                 | | |  |  |  VCLAMP
*                 | | |  |  |  | GND(REFERENCE)
.SUBCKT SMX10114  1 2 3A 4A 5    100
*
* DC PSRR FIX
J1 11 16 13 SMX10114QA
EPSRR- 16 2 TABLE {-V(4)} = (0,150U) (20,-50U)
J2 12 15 14 SMX10114QB
EPSRR+ 1 15 TABLE {V(3)} = (0,150U) (20,-50U)
*
* GMIN FIX
* GMIN = 1E-12, IF CHANGED MAKE RGI = -1/GMIN
RGS1 13 16 -1T
RGD1 16 11 -1T
RGS2 14 15 -1T
RGD2 12 15 -1T
*
RC1 4 11 1.67K
RC2 4 12 1.67K
C1 11 12 4.219P
RE1 13 10 667
RE2 14 10 667
GIEE 3 10 TABLE {V(3,4)} = (0,0) (2,0) (3,497U)
CE 10 100 12.59P
RE 10 100 402.4K
RP 3 4 8.564K
*
* CMRR FIX
GCM1 100 83 10 100 1
RCM1 83 84 1
LCM1 84 100 1.592U
GCM2 100 85 83 100 1
RCM2 85 86 1
LCM2 86 100 0.1592U
RCM3 86 100 10
GCM 100 21 85 100 52.15N
*
GA 21 100 11 12 598.8U
*
* PSRR VS FREQ FIX
GPSRR- 21 100 88 100 1
GVP- 100 88 4 100 1
RVP- 88 100 1
LVP- 88 100 0.1P
GPSRR+ 21 100 89 100 1
GVP+ 100 89 3 100 1
RVP+ 89 100 1
LVP+ 89 100 10P
*
R2 21 100 100K
C2 21 22 10P
GB 22 100 21 100 38.8
*
* VOLTAGE CLAMP
*RCL 9 100 100K
*VICL1 9 53
*VICL2 54 53
*RVOUT 54 55 10K
*EOUT 55 100 5 100 1
*WCL3 54 56 VICL3 CL
*RX 56 100 100K
*ICL+ 56 100 4M
*WCL4 54 57 VICL4 CL
*RY 57 100 100K
*ICL- 100 57 4M
*ECL1 47 100 9 100 1
*WCL1 47 48 VICL1 CL
*D8 48 49 SMX10114DD
*.MODEL SMX10114DD D (IS=1.075U)
*VICL3 49 6
*ECL2 52 100 9 100 1
*WCL2 52 51 VICL2 CL
*D9 50 51 SMX10114DE
*.MODEL SMX10114DE D (IS=15.28N)
*VICL4 6 50
*.MODEL CL ISWITCH (ION=2U IOFF=0 RON=1 ROFF=0.1MEG)
*
* END OF VCLAMP SECTION
RO2 22 100 31
D1 22 31 SMX10114DA
D2 31 22 SMX10114DC
EC 31 100 5 100 1.0
*
* I(VCC) FIX
RO1 22 6 19
VIOUT 6 5 0
D5 3 7 SMX10114DB
R5 7 100 1MEG
F5 7 100 VIOUT 1
D6 8 4 SMX10114DB
R6 8 100 1MEG
F6 8 100 VIOUT 1
*
* POWER OFF FIX
VIVP+ 3A 3
WVP+ 3 3B VIVP+ CL1
VIVP- 4 4A
WVP- 4 4B VIVP- CL1
.MODEL CL1 ISWITCH(
+        RON = 0.1
+       ROFF = 0.19MEG
+        ION = 0.5U
+       IOFF = 1N
+ )
*
* CLIPPING FIX
D3 5 24 SMX10114DB
EVC 3B 24 TABLE {V(3)} = (0,0.818) (5,2.258) (10,2.193) (15,2.268)
D4 25 5 SMX10114DB
EVE 25 4B TABLE {-V(4)} = (0,0.806) (5,2.186) (10,2.271) (15,2.286)
*
.MODEL SMX10114DA D (
+         IS = 13.11E-12
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL SMX10114DC D (
+         IS = 2.598E-6
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL SMX10114DB D (
+         IS = 0.8F
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL SMX10114QA PJF (
+        VTO = -1
+       BETA = 1M
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CGS = 0
+        CGD = 0
+         PB = 1
+         IS = 35E-12
+         KF = 0
+         AF = 1
+         FC = .5
+          N = 1
+        ISR = 0
+         NR = 2
+      ALPHA = 0
+         VK = 0
+          M = .5
+      VTOTC = 0
+    BETATCE = 0
+        XTI = 3
+ )
.MODEL SMX10114QB PJF (
+        VTO = -1.00116
+       BETA = 1M
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CGS = 0
+        CGD = 0
+         PB = 1
+         IS = 59.5E-12
+         KF = 0
+         AF = 1
+         FC = .5
+          N = 1
+        ISR = 0
+         NR = 2
+      ALPHA = 0
+         VK = 0
+          M = .5
+      VTOTC = 0
+    BETATCE = 0
+        XTI = 3
+ )
.ENDS SMX10114
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt TL082    1 2 3 4 5
*
  c1   11 12 2.412E-12
  c2    6  7 18.00E-12
  css  10 99 5.400E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 3.467E6 -1E3 1E3 3E6 -3E6
  ga    6  0 11 12 339.3E-6
  gcm   0  6 10 99 17.01E-9
  iss  10  4 dc 234.0E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   3 11 2.947E3
  rd2   3 12 2.947E3
  ro1   8  5 50
  ro2   7 99 170
  rp    3  4 20.00E3
  rss  10 99 854.7E3
  vb    9  0 dc 0
  vc    3 53 dc 1.500
  ve   54  4 dc 1.500
  vlim  7  8 dc 0
  vlp  91  0 dc 50
  vln   0 92 dc 50
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx NJF(Is=2.500E-12 Beta=984.2E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt TL084    1 2 3 4 5
*
  x_tl084 1 2 3 4 5 TL082
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt uA709    1 2 3 4 5 6 7
*
  c1   11 12 28.87E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 14.32E3 -1E3 1E3 10E3 -10E3
  ga    6  0 11 12 31.42E-3
  gcm   0  6 10 99 993.6E-9
  iee  10  4 dc 2.000E-3
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 31.83
  rc2   3 12 31.83
  re1  13 10 5.962
  re2  14 10 5.962
  ree  10 99 99.98E3
  ro1   8  5 50
  ro2   7 99 100
  rp    3  4 45.01E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 50
  vln   0 92 dc 50
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=5.000E3)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt ua709a   1 2 3 4 5 6 7
*
  c1   11 12 57.74E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 477.5E3 -1E3 1E3 480E3 -480E3
  ga    6  0 11 12 1.257E-3
  gcm   0  6 10 99 3.974E-9
  iee  10  4 dc 100.2E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 795.8
  rc2   3 12 795.8
  re1  13 10 277.9
  re2  14 10 277.9
  ree  10 99 1.996E6
  ro1   8  5 75
  ro2   7 99 75
  rp    3  4 12.50E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 100
  vln   0 92 dc 100
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=500)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |  compensation
*                | | | | | / \
.subckt ua709c   1 2 3 4 5 6 7
*
  c1   11 12 57.74E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 477.5E3 -1E3 1E3 480E3 -480E3
  ga    6  0 11 12 1.257E-3
  gcm   0  6 10 99 39.74E-9
  iee  10  4 dc 100.6E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 795.8
  rc2   3 12 795.8
  re1  13 10 276.8
  re2  14 10 276.8
  ree  10 99 1.988E6
  ro1   8  5 75
  ro2   7 99 75
  rp    3  4 11.69E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 100
  vln   0 92 dc 100
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=166.7)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt uA741    1 2 3 4 5
*
  c1   11 12 8.661E-12
  c2    6  7 30.00E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 10.61E6 -1E3 1E3 10E6 -10E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.836E3
  re2  14 10 1.836E3
  ree  10 99 13.19E6
  ro1   8  5 50
  ro2   7 99 100
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt ua771    1 2 3 4 5
*
  c1   11 12 3.750E-12
  c2    6  7 7.500E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 55.92E6 -1E3 1E3 56E6 -56E6
  ga    6  0 11 12 141.4E-6
  gcm   0  6 10 99 44.71E-9
  iss   3 10 dc 97.50E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   4 11 7.074E3
  rd2   4 12 7.074E3
  ro1   8  5 60
  ro2   7 99 40
  rp    3  4 10.00E-3
  rss  10 99 2.051E6
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx PJF(Is=25.00E-12 Beta=205.0E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt ua771a   1 2 3 4 5
*
  c1   11 12 3.750E-12
  c2    6  7 7.500E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 55.92E6 -1E3 1E3 56E6 -56E6
  ga    6  0 11 12 141.4E-6
  gcm   0  6 10 99 14.14E-9
  iss   3 10 dc 97.50E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   4 11 7.074E3
  rd2   4 12 7.074E3
  ro1   8  5 60
  ro2   7 99 40
  rp    3  4 10.00E-3
  rss  10 99 2.051E6
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx PJF(Is=25.00E-12 Beta=205.0E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt ua772    1 2 3 4 5
*
  c1   11 12 3.750E-12
  c2    6  7 7.500E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 29.82E6 -1E3 1E3 30E6 -30E6
  ga    6  0 11 12 141.4E-6
  gcm   0  6 10 99 44.71E-9
  iss   3 10 dc 97.50E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   4 11 7.074E3
  rd2   4 12 7.074E3
  ro1   8  5 75
  ro2   7 99 75
  rp    3  4 10.00E-3
  rss  10 99 2.051E6
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx PJF(Is=25.00E-12 Beta=205.0E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt ua772a   1 2 3 4 5
*
  c1   11 12 3.750E-12
  c2    6  7 7.500E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 55.92E6 -1E3 1E3 56E6 -56E6
  ga    6  0 11 12 141.4E-6
  gcm   0  6 10 99 14.14E-9
  iss   3 10 dc 97.50E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   4 11 7.074E3
  rd2   4 12 7.074E3
  ro1   8  5 60
  ro2   7 99 40
  rp    3  4 10.00E-3
  rss  10 99 2.051E6
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx PJF(Is=25.00E-12 Beta=205.0E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt ua772l   1 2 3 4 5
*
  c1   11 12 3.750E-12
  c2    6  7 7.500E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 55.92E6 -1E3 1E3 56E6 -56E6
  ga    6  0 11 12 141.4E-6
  gcm   0  6 10 99 44.71E-9
  iss   3 10 dc 97.50E-6
  hlim 90  0 vlim 1K
  j1   11  2 10 jx
  j2   12  1 10 jx
  r2    6  9 100.0E3
  rd1   4 11 7.074E3
  rd2   4 12 7.074E3
  ro1   8  5 60
  ro2   7 99 40
  rp    3  4 10.00E-3
  rss  10 99 2.051E6
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 25
  vln   0 92 dc 25
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model jx PJF(Is=25.00E-12 Beta=205.0E-6 Vto=-1)
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | output
*                | | | | |
.subckt ua798    1 2 3 4 5
*
  c1   11 12 8.660E-12
  c2    6  7 5.000E-12
  dc    5 53 dy
  de   54  5 dy
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2),(3,0),(4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 24.49E6 -1E3 1E3 24E6 -24E6
  ga    6  0 11 12 31.42E-6
  gcm   0  6 10 99 993.5E-12
  iee   3 10 dc 3.100E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   4 11 31.83E3
  rc2   4 12 31.83E3
  re1  13 10 14.12E3
  re2  14 10 14.12E3
  ree  10 99 64.52E6
  ro1   8  5 270
  ro2   7 99 260
  rp    3  4 15.02E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 70
  vln   0 92 dc 70
.model dx D(Is=800.0E-18)
.model dy D(Is=800.00E-18 Rs=1m Cjo=10p)
.model qx PNP(Is=800.0E-18 Bf=30)
.ends
*$
*-----------------------------------------------------------------------------

*** Voltage comparators

* The parameters in this comparator library were derived from data sheets for
* each parts.  The macromodel used was developed by MicroSim Corporation, and
* is produced by the "Parts" option to PSpice.
*
* Although we do not use it, another comparator macro model is described in:
*
*       An Integrated-Circuit Comparator Macromodel
*         by Ian Getreu, Andreas Hadiwidjaja, and Johan Brinch
*       IEEE Journal of Solid-State Circuits, Vol. SC-11, no. 6, Dec. 1976
*
* This reference covers the considerations that go into duplicating the
* behavior of voltage comparators.
*
* The comparators are modelled at room temperature.  The macro model does not
* track changes with temperature.  This library file contains models for
* nominal, not worst case, devices.
*$
*
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | | output ground
*                | | | | | |
.subckt LM111    1 2 3 4 5 6
*
  f1    9  3 v1 1
  iee   3  7 dc 100.0E-6
  vi1  21  1 dc .45
  vi2  22  2 dc .45
  q1    9 21  7 qin
  q2    8 22  7 qin
  q3    9  8  4 qmo
  q4    8  8  4 qmi
.model qin PNP(Is=800.0E-18 Bf=833.3)
.model qmi NPN(Is=800.0E-18 Bf=1002)
.model qmo NPN(Is=800.0E-18 Bf=1000 Cjc=1E-15 Tr=118.8E-9)
  e1   10  6  9  4  1
  v1   10 11 dc 0
  q5    5 11  6 qoc
.model qoc NPN(Is=800.0E-18 Bf=34.49E3 Cjc=1E-15 Tf=364.6E-12 Tr=79.34E-9)
  dp    4  3 dx
  rp    3  4 6.122E3
.model dx  D(Is=800.0E-18 Rs=1)
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | | output ground
*                | | | | | |
.subckt LM119    1 2 3 4 5 6
*
  f1    3  9 v1 1
  iee   7  4 dc 100.0E-6
  q1    9  2  7 qin
  q2    8  1  7 qin
  q3    9  8  3 qmo
  q4    8  8  3 qmi
.model qin NPN(Is=800.0E-18 Bf=333.3)
.model qmi PNP(Is=800.0E-18 Bf=1002)
.model qmo PNP(Is=800.0E-18 Bf=1000 Cjc=1E-15 Tr=59.42E-9)
  e1   10  6  3  9  1
  v1   10 11 dc 0
  q5    5 11  6 qoc
.model qoc NPN(Is=800.0E-18 Bf=41.38E3 Cjc=1E-15 Tf=23.91E-12 Tr=24.01E-9)
  dp    4  3 dx
  rp    3  4 5.556E3
.model dx  D(Is=800.0E-18 Rs=1)
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | |
.subckt LM139    1 2 3 4 5
*
  f1    9  3 v1 1
  iee   3  7 dc 100.0E-6
  vi1  21  1 dc .75
  vi2  22  2 dc .75
  q1    9 21  7 qin
  q2    8 22  7 qin
  q3    9  8  4 qmo
  q4    8  8  4 qmi
.model qin PNP(Is=800.0E-18 Bf=2.000E3)
.model qmi NPN(Is=800.0E-18 Bf=1002)
.model qmo NPN(Is=800.0E-18 Bf=1000 Cjc=1E-15 Tr=475.4E-9)
  e1   10  4  9  4  1
  v1   10 11 dc 0
  q5    5 11  4 qoc
.model qoc NPN(Is=800.0E-18 Bf=20.69E3 Cjc=1E-15 Tf=3.540E-9 Tr=472.8E-9)
  dp    4  3 dx
  rp    3  4 37.50E3
.model dx  D(Is=800.0E-18 Rs=1)
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | |
.subckt LM193    1 2 3 4 5
*
  x_lm193 1 2 3 4 5 LM139
*
* the LM193 is identical to the LM139, but in a different package
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | | output ground
*                | | | | | |
.subckt LM211    1 2 3 4 5 6
*
  x_lm211 1 2 3 4 5 6 LM111
*
* the LM211 is identical to the LM111, but has a more limited temp. range
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | | output ground
*                | | | | | |
.subckt LM219    1 2 3 4 5 6
*
  x_lm219 1 2 3 4 5 6 LM119
*
* the LM219 is identical to the LM119, but has a more limited temp. range
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | |
.subckt LM239    1 2 3 4 5
*
  x_lm239 1 2 3 4 5 LM139
*
* the LM239 is identical to the LM139, but has a more limited temp. range
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | |
.subckt LM293    1 2 3 4 5
*
  x_lm293 1 2 3 4 5 LM139
*
* the LM293 is identical to the LM239, but in a different package
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | | output ground
*                | | | | | |
.subckt LM311    1 2 3 4 5 6
*
f1    9  3 v1 1
iee   3  7 dc 100.0E-6
vi1  21  1 dc .45
vi2  22  2 dc .45
q1    9 21  7 qin
q2    8 22  7 qin
q3    9  8  4 qmo
q4    8  8  4 qmi
.model qin PNP(Is=800.0E-18 Bf=500)
.model qmi NPN(Is=800.0E-18 Bf=1002)
.model qmo NPN(Is=800.0E-18 Bf=1000 Cjc=1E-15 Tr=124.2E-9)
e1   10  6  9  4  1
v1   10 11 dc 0
q5    5 11  6 qoc
.model qoc NPN(Is=800.0E-18 Bf=206.9E3 Cjc=1E-15 Tf=7.855E-12 Tr=83.83E-9)
dp    4  3 dx
rp    3  4 7.087E3
.model dx  D(Is=800.0E-18)
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | | output ground
*                | | | | | |
.subckt LM319    1 2 3 4 5 6
*
  x_lm319 1 2 3 4 5 6 LM119
*
* the LM319 is identical to the LM119, but has a more limited temp. range
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | |
.subckt LM339    1 2 3 4 5
*
  x_lm339 1 2 3 4 5 LM139
*
* the LM339 is identical to the LM139, but has a more limited temp. range
*
.ends
*$
*
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | |
.subckt LM393    1 2 3 4 5
*
  x_lm393 1 2 3 4 5 LM139
*
* the LM393 is identical to the LM339, but in a different package
*
.ends
*$
*-----------------------------------------------------------------------------
* connections:   non-inverting input
*                | inverting input
*                | | positive power supply
*                | | | negative power supply
*                | | | | open collector output
*                | | | | |
.subckt LM3302   1 2 3 4 5
*
  x_lm3302 1 2 3 4 5 LM139
*
* the LM3302 is identical to the LM139, but has a more limited temp. range
*
.ends
*$
*-----------------------------------------------------------------------------

*** Voltage regulators (positive)

.SUBCKT x_LM78XX Input Output Ground PARAMS:
+       Av_feedback=1665, R1_Value=1020
*
* SERIES 3-TERMINAL POSITIVE REGULATOR
*
* Note: This regulator is based on the LM78XX series of
*       regulators (also the LM140 and LM340).  The model
*       will cause some current to flow to Node 0 which
*       is not part of the actual voltage regulator circuit.
*
* Band-gap voltage source:
*
*       The source is off when Vin<3V and fully on when Vin>3.7V.
*       Line regulation and ripple rejection) are set with
*       Rreg= 0.5 * dVin/dVbg.  The temperature dependence of this
*       circuit is a quadratic fit to the following points:
*
*                                T         Vbg(T)/Vbg(nom)
*                               ---        ---------------
*                                0            .999
*                               37.5            1
*                               125           .990
*
*       The temperature coefficient of Rbg is set to 2 * the band gap
*       temperature coefficient.  Tnom is assumed to be 27 deg. C and
*       Vnom is 3.7V
*
Vbg 100 0 DC 7.4V
Sbg (100,101),(Input,Ground) Sbg1
Rbg 101 0 1 TC=1.612E-5,-2.255E-6
Ebg (102,0),(Input,Ground) 1
Rreg 102 101 7k
.MODEL Sbg1 VSWITCH (Ron=1 Roff=1MEG Von=3.7 Voff=3)
*
* Feedback stage
*
*       Diodes D1,D2 limit the excursion of the amplifier
*       outputs to being near the rails.  Rfb, Cfb Set the
*       corner frequency for roll-off of ripple rejection.

*
*       The opamp gain is given by:  Av = (Fores/Freg) * (Vout/Vbg)
*       where Fores = output impedance corner frequency
*                     with Cl=0 (typical value about 1MHz)
*             Freg  = corner frequency in ripple rejection
*                     (typical value about 600 Hz)
*             Vout  = regulator output voltage (5,12,15V)
*             Vbg   = bandgap voltage (3.7V)
*
*       Note: Av is constant for all output voltages, but the
*       feedback factor changes. If Av=2250, then the
*       Av*Feedback factor is as given below:
*
*                                 Vout     Av*Feedback factor
*                                 ----     ------------------
*                                   5          1665
*                                  12           694
*                                  15           550
*
Rfb 9 8 1MEG
Cfb 8 Ground 265PF
Eopamp 105 0 VALUE={2250*v(101,0)+Av_feedback*v(Ground,8)}
Vgainf 200 0 {Av_feedback}
Rgainf 200 0 1
*Eopamp 105 0 POLY(3),(101,0),(Ground,8),(200,0) 0 2250 0 0 0 0 0 0 1
Ro 105 106 1k
D1 106 108 Dlim
D2 107 106 Dlim
.MODEL Dlim D (Vj=0.7)
Vl1 102 108 DC 1
Vl2 107 0 DC 1
*
* Quiescent current modelling
*
*       Quiescent current is set by Gq, which draws a current
*       proportional to the voltage drop across the regulator and
*       R1 (temperature coefficient .1%/deg C).  R1 must change
*       with output voltage as follows:  R1 = R1(5v) * Vout/5v.
*
Gq (Input,Ground),(Input,9) 2.0E-5
R1 9 Ground {R1_Value} TC=0.001
*
* Output Stage
*
*       Rout is used to set both the low frequency output impedence
*       and the load regulation.
*
Q1 Input 5 6 Npn1
Q2 Input 6 7 Npn1 10
.MODEL Npn1 NPN (Bf=50 Is=1E-14)
* Efb Input 4 VALUE={v(Input,Ground)+v(0,106)}
Efb Input 4 POLY(2),(Input,Ground),(0,106) 0 1 1
Rb 4 5 1k TC=0.003
Re 6 7 2k
Rsc 7 9 0.275 TC=1.136E-3,-7.806E-6
Rout 9 Output 0.008
*
* Current Limit
*
Rbcl 7 55 290
Qcl 5 55 9 Npn1
Rcldz 56 55 10k
Dz1 56 Input Dz
.MODEL Dz D (Is=0.05p Rs=3 Bv=7.11 Ibv=0.05u)
.ENDS
*$
*
*---------------------------------------------------------------LM7805C
.SUBCKT LM7805C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
*---------------------------------------------------------------uA7805C
.SUBCKT UA7805C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
* MANUFACTURERS PART NO.= UA7805  (TEXAS INTERNATIONAL)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMP. DEPENDENT MODEL OF THE UA7805
* REGULATOR.
*
*------------------------------------------------------------------------------
*
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT.  IT
* INCLUDES POWER-UP AND POWER-DOWN EFFECTS.
* IT MAY BE NECESSARY TO SET ITL1=300 ITL2=300 WITH THE .OPTIONS COMMAND
* FOR CONVERGENCE.  THESE SETTINGS DETERMINE THE NUMBER OF ITERATIONS
* ALLOWED FOR THE CALCULATION OF THE DC AND BIAS PT VALUES WHEN THE
* STARTING POINT IS  CONSIDERED "BLIND" OR AN "EDUCATED GUESS".
* OTHER SETTINGS MAY WORK, BUT HAVE NOT BEEN TESTED YET.
*
*
*
.SUBCKT UA7805/TEMP  1  2   3
*                    |  |   |
*                   IN  |   |
*                      OUT  |
*                          GND
*




*** VOLTAGE REFERENCE AND BIAS CURRENT SECTION ***
DZ1  4 1 DZ1
.MODEL DZ1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.5
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -0.001481
+       TBV2 = -1.85167E-5
+       TRS1 = 0
+       TRS2 = 0
+ )
RQ   4 17 112090 TC=0.003483, -4.9343E-6
RR   17 18 4.7 TC=0.003449, -5.495E-6
DR   16 18 DR
.MODEL DR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.2651
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 1.805303E-4
+       TBV2 = -2.461378E-6
+       TRS1 = 0
+       TRS2 = 0
+ )
RZ 16 18 1MEG
L1 16 3 IND1 0.796M
.MODEL IND1 IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 0.00236
+        TC2 = 1.24436E-5
+ )
*** ERROR AMPLIFIER SECTION ***
EP 22 3 17 15 300
RO 22 6 25
DC- 3 6 DCLAMP
DC+ 6 19 DCLAMP
.MODEL DCLAMP D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
V+ 19 23 DC -1
E+ 23 3 1 3 1
RP 6 7 50
CPZ 7 3 0.5U
*** QUIESCENT CURRENT ***
GB 1 9 17 3 0.5002M
RQUIES 12 3 3396 TC=0.006886, 4.655264E-5
*** SHORT CIRCUIT AND FOLDBACK CURRENT ***
DBL 9 8 DBL
.MODEL DBL D(
+         IS = 1E-4
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
EB 8 3 7 3 2
RC 1 14 0.2
DC 14 13 DC
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1.617
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
RB 9 11 100
QP 13 11 5 QP
.MODEL QP NPN(
+         IS = 1E-12
+         BF = 70K
+         NF = 1
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
DCL 9 10 DCL
.MODEL DCL D(
+         IS = 1E-4
+         RS = 0
+          N = 2
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
QCL 10 20 12 QLIMIT
.MODEL QLIMIT NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
RSC 5 12 .5076
RBCL 20 5 1600
RFBCL 1 21 51.17K TC= 0.002528, -1.5164E-5
DZFB 20 21 DZFB
.MODEL DZFB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 15.26
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -9.5474743E-4
+       TBV2 = 1.478994E-5
+       TRS1 = 0
+       TRS2 = 0
+ )
R24 15 3 600
R23 12 15 1850
*** OUTPUT RESISTANCE ***
ROUT 12 2 0.036 TC=0.002616, -1.50463E-5
DDIS 12 1 DMOD
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 0.7
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS UA7805/TEMP
*$
*
*
* GENERIC FUNCTIONAL EQUIVALENT = DT831031B
* TYPE: DIODE
* SUBTYPE: VOLTAGE_REF_TC

* THIS FILE CONTAINS 5 MODELS AT VARIOUS TEST CONDITIONS.
* PARAMETER MODELS EXTRACTED FROM MEASURED DATA

* RAD: PRERAD
* TEMP= 27

*** CAUTION: MODEL IS VALID FOR OPERATION IN THE REVERSE REGION ONLY!

.SUBCKT DT831031B/27C  99  2
D1  2   99   DLEAK
R1  2   99   1E12
V2  5   99   20.73
D2  2   5   DBLOCK
C1  2   99   5.5E-11
.MODEL DLEAK    D       (
+         IS = 3.219715E-12
+         RS = 0.0609964
+          N = 58.2632139
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL DBLOCK   D       (
+         IS = 3.066643E-11
+         RS = 1.6578749
+          N = 8.1826239
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.ENDS
*$
*
* RAD: PRERAD
* TEMP= -55

*** CAUTION: MODEL IS VALID FOR OPERATION IN THE REVERSE REGION ONLY!

.SUBCKT DT831031B/-55C  99  2
D1  2   99   DLEAK
R1  2   99   1E12
V2  5   99   20.93
D2  2   5   DBLOCK
C1  2   99   4.65E-11
.MODEL DLEAK    D       (
+         IS = 2.294595E-14
+         RS = 0.0609964
+          N = 62.9736183
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL DBLOCK   D       (
+         IS = 2.03286E-11
+         RS = 1.7841132
+          N = 9.602096
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.ENDS
*$
*
* RAD: PRERAD
* TEMP= 125

*** CAUTION: MODEL IS VALID FOR OPERATION IN THE REVERSE REGION ONLY!

.SUBCKT DT831031B/125C  99  2
D1  2   99   DLEAK
R1  2   99   1E12
V2  5   99   20.14
D2  2   5   DBLOCK
C1  2   99   6.8E-11
.MODEL DLEAK    D       (
+         IS = 1.569829E-12
+         RS = 0.0609964
+          N = 39.3712792
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL DBLOCK   D       (
+         IS = 1.612864E-11
+         RS = 2.4440014
+          N = 7.4242884
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.ENDS
*$
*
* TYPE: DIODE
* SUBTYPE: VOLTAGE_REF_TC

* THE FOLLOWING SECTION CONTAINS 2 PARAMETER SETS AT VARIOUS POST NEUTRON
* RADIATION LEVELS.
* PARAMETER SETS EXTRACTED FROM MEASURED DATA.

*** CAUTION: MODEL IS VALID FOR OPERATION IN THE REVERSE REGION ONLY!
*** CAUTION: USE ONLY AT TEMPERATURE SPECIFIED.  ANY DEVIATION FROM THIS
***          TEMPERATURE WILL PRODUCE INCORRECT RESULTS.

* RAD: 2.2E13
* TYPE: NEUTRON
* TEMP: 27
*
.SUBCKT DT831031B/27C/RAD1  99  2
D1  2   99   DLEAK
R1  2   99   1E12
V2  5   99   20.71
D2  2   5   DBLOCK
C1  2   99   6E-11
.MODEL DLEAK    D       (
+         IS = 3.258506E-10
+         RS = 15.2165394
+          N = 80.8147666
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL DBLOCK   D       (
+         IS = 3.80381E-11
+         RS = 1.438611
+          N = 8.32254
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.ENDS
*$
*
* RAD: 2.73E14
* TYPE: NEUTRON
* TEMP: 27
*
.SUBCKT DT831031B/27C/RAD2  99  2
D1  2   99   DLEAK
R1  2   99   1E12
V2  5   99   20.40
D2  2   5   DBLOCK
C1  2   99   4.7E-11
.MODEL DLEAK    D       (
+         IS = 1.772633E-10
+         RS = 0.0609964
+          N = 68.8487735
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL DBLOCK   D       (
+         IS = 8.377173E-12
+         RS = 2.2593796
+          N = 8.2245024
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.ENDS
*$
*
* MANUFACTURERS PART NO. = L161AL  (SILICONIX)
* SUBTYPE: COMPARATOR
* THIS IS A PRE-RAD MODEL AT 27 C OF THE L161AL
* THIS MODEL MAY BE USED FOR ALL OF THE FOLLOWING DEVICES :
* L161AP
* L161AL
*
*
** THE FOLLOWING ARE THE LIMITATIONS OF THIS MODEL:
*
* THIS MODEL IS A TRANSISTOR LEVEL MODEL OF THE SILICONIX L161 VOLTAGE
* COMPARATOR WHICH FOLLOWS THE SCHEMATIC FROM THE DATA SHEET AND THE
* PRODUCT  SPEC.  THIS MODEL DOES NOT SIMULATE VOS AND IOS.  IT DOES
* SIMULATE IBT, VOL,  VOH, AND IS ACCORDING TO PRODUCT SPEC LIMITS.  THE
* MODEL SIMULATES +SR  WITHIN 5% OF THE SILICONIX DATA SHEET VALUES(PAGE 8-
* 46).  IT DOES NOT  SIMULATE -SR.  -SR FOR THE ACTUAL DEVICE IS APPROXIMATELY
* 3 TIMES FASTER  THAN THE MODEL SIMULATION.  THE MODEL SIMULATES
* RESPONSE TIME (TRLH) FOR  A 100MV OVERDRIVE WITHIN 12% OF THE SILICONIX
* DATA SHEET(PAGE 8-47) AND  TRHL WITHIN 20%.  IT DOES NOT SIMULATE RESPONSE
* TIME FOR A 5MV OVERDRIVE.
* THE ACTUAL DEVICE IS 2.5 TIMES FASTER FOR TRLH AND IS 5 TIMES FASTER FOR
* TRHL.  THE MODEL DOES NOT SIMULATE A 20MV OVERDRIVE.  THE ACTUAL DEVICE
* IS 1.3 TIMES FASTER FOR TRLH AND 2.3 FASTER FOR TRHL.
*
*  CONNECTIONS:   NON-INVERTING INPUT
*                 |  INVERTING INPUT
*                 |  |  POSITIVE POWER SUPPLY
*                 |  |  |  NEGATIVE POWER SUPPLY
*                 |  |  |  |  OUTPUT
*                 |  |  |  |  |  ISET
*                 |  |  |  |  |  |
.SUBCKT L161      9  7  1  8  10 14
*
Q1 8 7 3 PNPNOM
QD1 4 4 8 NPNNOM
Q2 8 9 6 PNPNOM
Q3A 3 3 2 PNPNOM
Q3B 4 3 2 PNPNOM 7
Q4A 6 6 2 PNPNOM
Q4B 5 6 2 PNPNOM 7
Q5 5 4 8 NPNNOM
Q6A 11 11 1 PNPNOM
Q6B 10 11 1 PNPNOM 2
Q6C 2 11 1 PNPNOM 2
Q7 10 5 8 NPNNOM 2
Q8 11 12 8 NPNNOM
Q9 1 13 12 NPNNOM
Q10 13 12 8 NPNNOM
J11 14 8 13 JNOM
.MODEL NPNNOM NPN  (
+         IS = 1.66E-16
+         BF = 100
+         NF = 1
+        VAF = 200
+        IKF = 7E-3
+        ISE = 0
+         NE = 1.5
+         BR = 1.1
+         NR = 1
+        VAR = 26
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 150
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 3
+         RC = 800
+        CJE = 1.35E-12
+        VJE = 0.964
+        MJE = 0.5
+         TF = 1E-9
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 1.35E-12
+        VJC = 0.663
+        MJC = 0.5
+       XCJC = 1
+         TR = 100E-9
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 1E-12
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL PNPNOM PNP  (
+         IS = 2.83E-17
+         BF = 40
+         NF = 1
+        VAF = 80
+        IKF = 0.1E-3
+        ISE = 0
+         NE = 1.5
+         BR = 4
+         NR = 1
+        VAR = 40
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 400
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 20
+         RC = 1400
+        CJE = 0.85E-12
+        VJE = 0.663
+        MJE = 0.5
+         TF = 100E-9
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 1.18E-12
+        VJC = 0.663
+        MJC = 0.5
+       XCJC = 1
+         TR = 100E-9
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 1E-12
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL JNOM NJF(
+        VTO = -18
+       BETA = 1E-5
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CGS = 0
+        CGD = 0
+         PB = 1
+         IS = 1E-14
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.ENDS L161
*$
*
*---------------------------------------------------------------LAS1505
.SUBCKT LAS1505 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
* MANUFACTURERS PART NO. = LM129AH/883B  (NATIONAL SEMICONDUCTOR)  
* TYPE: IC_LINEAR  
* SUBTYPE: REFERENCE  
* THIS FILE CONTAINS 1 PRERAD TEMPERATURE DEPENDENT MACROMODEL OF THE LM129AH  
* VOLTAGE REFERENCE  
* CREATION DATE :  9-24-92  
*  
* PLEASE NOTE THE FOLLOWING:  
*  
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT.  
* IT NEEDS TO BE RUN WITH VERSION 4.03 OR HIGHER OF PSPICE DUE TO THE  
* TEMPERATURE COEFFICIENTS IN THE MODEL FOR THE INDUCTORS AND THE DIODE  
* BREAKDOWN VOLTAGE.  IT IS NECESSARY TO SET ITL1=300 ITL2=300 WITH THE  
* .OPTIONS COMMAND FOR 100% CONVERGENCE.  THESE SETTINGS DETERMINE THE  
* NUMBER OF ITERATIONS ALLOWED FOR THE CALCULATION OF THE DC AND BIAS PT  
* VALUES WHEN THE STARTING POINT IS CONSIDERED "BLIND" OR AN "EDUCATED GUESS".  
* OTHER SETTINGS MAY WORK, BUT HAVE NOT BEEN TESTED YET.  
*  
*------------------------------------------------------------------------------  
*  
*  
.SUBCKT LM129  1   2  
**********     |   |  
*********      + (CATHODE)  
***********        - (ANODE)  
*  
DR 3 1 DMOD  
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 6.847
+        IBV = .001
+ )
CR 3 1 CR 300PF  
.MODEL CR CAP(
*PSPICE (MicroSim) Specific Parameters Follow
+          C = 1
+        VC1 = 0
+        VC2 = 0
+        TC1 = 0.44
+        TC2 = 0.0055
+ )
RDR 3 4 0.6211 TC=2.7447E-4, 1.2663E-5  
LDR 4 2 LDR 0.0247MH  
.MODEL LDR IND(
*PSPICE (MicroSim) Specific Parameters Follow
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 8.5774E-3
+        TC2 = 2.4348E-5
+ )
RLDR 4 2 50  
.ENDS LM129  
*$
*  
* RAD: PRERAD  
*  
* TEMP= -55  
*  
*** NOTE: TRR MEASUREMENT WAS MADE @ 10MA/10MA/2.5MA  
*  
*** CAUTION: THE MEASURED TRR AND THE PSPICE CKT. SIMULATED TRR ARE DIFFERENT  
*            THIS COULD POTENTIALLY LEAD TO ERRORS IN CKT. SIMULATIONS IF USED  
*            AS A RECTIFIER OR SWITCHING DIODE  
*  
* MEASURED TRR = 627.0NS, SIMULATED TRR = 493.0NS.  
*  
.SUBCKT LM129/-55C  99  2  
D1  2   99   DLEAK1  
R1  2   99   1E12  
R2  6   99   0.81  
M1  2   2   6   8   MOS1  
R3  6   8   1E12  
V2  10  99   5.45  
D2  2   10  DLEAK2  
D3  99   2   DFOR  
.MODEL DLEAK1   D       (
+         IS = 2.76E-16
+         RS = 0.6745712
+          N = 14.579
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL MOS1     NMOS    (
+      LEVEL = 1
+        VTO = 6.802
+         KP = 1E7
+      GAMMA = 0
+        PHI = .6
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CBD = 0
+        CBS = 0
+         IS = 1E-14
+         PB = .8
+       CGSO = 0
+       CGDO = 0
+       CGBO = 0
+        RSH = 0
+         CJ = 0
+         MJ = .5
+       CJSW = 0
+       MJSW = .33
+         JS = 1E-08
+        TOX = .0000001
+        NSS = 0
+        NFS = 0
+        TPG = 1
+         XJ = 0
+         LD = 0
+         UO = 600
+      UCRIT = 10000
+       UEXP = 0
+       UTRA = 0
+       VMAX = 0
+       NEFF = 1
+        XQC = 1
+         KF = 0
+         AF = 1
+         FC = .5
+      DELTA = 0
+      THETA = 0
+        ETA = 0
+      KAPPA = .2
+ )
.MODEL DLEAK2   D       (
+         IS = 5E-13
+         RS = 2E3
+          N = 1.1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL DFOR     D       (
+         IS = 1.237167E-10
+         RS = 21.0306341
+          N = 1.5903301
+         TT = 6.80E-7
+        CJO = 2.216063E-11
+         VJ = 0.7379787
+          M = 0.2379013
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = 0.5
+         BV = 1E5
+        IBV = .001
+ )
.ENDS LM129/-55C
*
*$
* RAD: PRERAD  
*  
* TEMP= 125  
*  
*** NOTE: TRR MEASUREMENT WAS MADE @ 10MA/10MA/2.5MA  
*  
*** CAUTION: THE MEASURED TRR AND THE PSPICE CKT. SIMULATED TRR ARE DIFFERENT  
*            THIS COULD POTENTIALLY LEAD TO ERRORS IN CKT. SIMULATIONS IF USED  
*            AS A RECTIFIER OR SWITCHING DIODE  
*  
* MEASURED TRR = 2.117US, SIMULATED TRR = 905.8NS.  
*  
.SUBCKT LM129/125C  99  2  
D1  2   99   DLEAK1  
R1  2   99   5E8  
R2  6   99   0.58  
M1  2   2   6   8   MOS1  
R3  6   8   1E15  
V2  10  99   6  
D2  2   10  DLEAK2  
D3  99   2   DFOR  
.MODEL DLEAK1   D       (
+         IS = 3E-14
+         RS = 0.6746
+          N = 11
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL MOS1     NMOS    (
+      LEVEL = 1
+        VTO = 6.984
+         KP = 1E7
+      GAMMA = 0
+        PHI = .6
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CBD = 0
+        CBS = 0
+         IS = 1E-18
+         PB = .8
+       CGSO = 0
+       CGDO = 0
+       CGBO = 0
+        RSH = 0
+         CJ = 0
+         MJ = .5
+       CJSW = 0
+       MJSW = .33
+         JS = 1E-08
+        TOX = .0000001
+        NSS = 0
+        NFS = 0
+        TPG = 1
+         XJ = 0
+         LD = 0
+         UO = 600
+      UCRIT = 10000
+       UEXP = 0
+       UTRA = 0
+       VMAX = 0
+       NEFF = 1
+        XQC = 1
+         KF = 0
+         AF = 1
+         FC = .5
+      DELTA = 0
+      THETA = 0
+        ETA = 0
+      KAPPA = .2
+ )
.MODEL DLEAK2   D       (
+         IS = 1E-12
+         RS = 2.3E3
+          N = 1.64
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL DFOR     D       (
+         IS = 1.5E-13
+         RS = 18
+          N = 1.05
+         TT = 1.2E-6
+        CJO = 2.88E-11
+         VJ = 0.35
+          M = 0.297
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = 0.860
+         BV = 1E5
+        IBV = .001
+ )
.ENDS LM129/125C
*$
* MANUFACTURERS PART NO. = LM129AH/883B  (NATIONAL SEMICONDUCTOR)  
* TYPE: IC_LINEAR  
* SUBTYPE: REFERENCE  
* THIS FILE CONTAINS 3 PRERAD SPICE2G.6 MACROMODELS AT 27 C, -55 C AND 125 C.  
* TEMPERATURE PARAMETER MODELS EXTRACTED FROM MEASURED DATA.  
* CREATION DATE : 07-05-90  
*  
*  
**************************************************************************  
* THE FOLLOWING MACROMODELS ARE SPICE2G.6 COMPATIBLE AND ARE FOR USE ONLY  
* AT THE TEMPERATURE INDICATED  
*  
* RAD: PRERAD  
*  
* TEMP= 27  
*  
*** NOTE: TRR MEASUREMENT WAS MADE @ 10MA/10MA/2.5MA  
*  
*** CAUTION: THE MEASURED TRR AND THE PSPICE CKT. SIMULATED TRR ARE DIFFERENT  
*            THIS COULD POTENTIALLY LEAD TO ERRORS IN CKT. SIMULATIONS IF USED  
*            AS A RECTIFIER OR SWITCHING DIODE  
*  
* MEASURED TRR = 1.305US, SIMULATED TRR = 544.4NS.  
*  
.SUBCKT LM129/27C  99  2  
D1  2   99   DLEAK1  
R1  2   99   9.99E11  
R2  6   99   0.6  
M1  2   2   6   8   MOS1  
R3  6   8   1E12  
V2  10  99   5.8  
D2  2   10  DLEAK2  
D3  99   2   DFOR  
.MODEL DLEAK1   D       (
+         IS = 1.66E-15
+         RS = 15.7046607
+          N = 12.12
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL MOS1     NMOS    (
+      LEVEL = 1
+        VTO = 6.885
+         KP = 1E7
+      GAMMA = 0
+        PHI = .6
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CBD = 0
+        CBS = 0
+         IS = 1E-14
+         PB = .8
+       CGSO = 0
+       CGDO = 0
+       CGBO = 0
+        RSH = 0
+         CJ = 0
+         MJ = .5
+       CJSW = 0
+       MJSW = .33
+         JS = 1E-08
+        TOX = .0000001
+        NSS = 0
+        NFS = 0
+        TPG = 1
+         XJ = 0
+         LD = 0
+         UO = 600
+      UCRIT = 10000
+       UEXP = 0
+       UTRA = 0
+       VMAX = 0
+       NEFF = 1
+        XQC = 1
+         KF = 0
+         AF = 1
+         FC = .5
+      DELTA = 0
+      THETA = 0
+        ETA = 0
+      KAPPA = .2
+ )
.MODEL DLEAK2   D       (
+         IS = 1.2E-16
+         RS = 2.2E3
+          N = 0.75
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL DFOR     D       (
+         IS = 4.16979E-10
+         RS = 8.541917
+          N = 1.6705528
+         TT = 7.4E-7
+        CJO = 2.724589E-11
+         VJ = 0.6060786
+          M = 0.2493594
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = 0.5
+         BV = 1E5
+        IBV = .001
+ )
.ENDS LM129/27C
*
*$
* MANUFACTURERS PART NO. = LM185BYH/883  (NATIONAL SEMICONDUCTOR)  
* TYPE: IC_LINEAR  
* SUBTYPE: REFERENCE  
* THIS FILE CONTAINS 3 PRE-RAD SPICE2G.6 COMPATIBLE MODELS AT VARIOUS TEMPS  
* OF THE LM185 TWO TERMINAL 1.2V REF.  
* PARAMETER MODELS EXTRACTED FROM MEASURED DATA  
* CREATION DATE : 07-02-90  
*  
*****CAUTION: THESE MODELS ARE ONLY GOOD FOR THE TEMPERATURE THEY WERE  
*             DEVELOPED AT.  
*  
* RAD: PRERAD  
* TEMP= 27  
*  
*** NOTE: TRR MEASUREMENT WAS MADE @ 10MA/10MA/2.5MA  
*  
*** CAUTION: THE MEASURED TRR AND THE PSPICE CKT. SIMULATED TRR ARE DIFFERENT  
*            THIS COULD POTENTIALLY LEAD TO ERRORS IN CKT. SIMULATIONS IF USED  
*            AS A RECTIFIER OR IN SWITCHING APPLICATIONS.  
*  
* MEASURED TRR = 1.03US, SIMULATED TRR = 720.4NS.  
*  
*  
.SUBCKT LM185/27C  99  2  
D1  2   99   DLEAK  
R1  2   99   1E12  
R2  6   99   0.12  
M1  2   2   6   8   MOS1  
R3  6   8   1E12  
D2  99   2   DFOR  
.MODEL DLEAK    D       (
+         IS = 2E-6
+         RS = 34.8744396
+          N = 53
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL MOS1     NMOS    (
+      LEVEL = 1
+        VTO = 2.512
+         KP = 1E7
+      GAMMA = 0
+        PHI = .6
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CBD = 0
+        CBS = 0
+         IS = 1E-14
+         PB = .8
+       CGSO = 0
+       CGDO = 0
+       CGBO = 0
+        RSH = 0
+         CJ = 0
+         MJ = .5
+       CJSW = 0
+       MJSW = .33
+         JS = 1E-08
+        TOX = .0000001
+        NSS = 0
+        NFS = 0
+        TPG = 1
+         XJ = 0
+         LD = 0
+         UO = 600
+      UCRIT = 10000
+       UEXP = 0
+       UTRA = 0
+       VMAX = 0
+       NEFF = 1
+        XQC = 1
+         KF = 0
+         AF = 1
+         FC = .5
+      DELTA = 0
+      THETA = 0
+        ETA = 0
+      KAPPA = .2
+ )
.MODEL DFOR     D       (
+         IS = 5.173495E-9
+         RS = 13.7420803
+          N = 2.0242147
+         TT = 9.74E-7
+        CJO = 7.094324E-11
+         VJ = 0.6122206
+          M = 0.2691849
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = 0.5
 +         BV = 1E5
+        IBV = .001
+ )
.ENDS LM185/27C
* 
*$
* MANUFACTURERS PART NO. = LM185BYH/883  (NATIONAL SEMICONDUCTOR)  
* TYPE: IC_LINEAR  
* SUBTYPE: REFERENCE  
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT SPICE2G.6 COMPATIBLE  
* MODEL OF THE LM185BYH ADJUSTABLE 1.2-5.3V REF  
* CREATION DATE : 11-28-90  
*  
*  
* LM185 ADJUSTABLE VOLTAGE REFERENCE "MACROMODEL" SUBCIRCUIT  
* THIS IS A TRANSISTOR LEVEL MODEL WHICH USES DEFAULT TRANSISTOR VALUES  
* (EBER'S MOLL) AND FOLLOWS THE SCHEMATIC OF THE NATIONAL DATA SHEET.  Q10  
* (ONE OF THE NPN TRANSISTORS IN THE BANDGAP REFERENCE SECTION) HAS A SCALING  
* FACTOR OF 10. THIS MODEL CAN BE USED WITH A .TEMP CARD.  IT ACCURATELY  
* SIMULATES CHANGE IN VREF WITH CHANGE IN CURRENT, ZOUT, AND IFEEDBACK.  
*  
***** CAUTION: THE MODEL EXCEEDS THE PRODUCT SPEC LIMIT FOR VREF AT 25 C BY  
*              2 MV AND AT 125 C BY 27 MV FOR IR = 8 UA AND IR = 100 UA.  
*  
* SINCE THIS IS A TRANSISTOR LEVEL MODEL(WITH 13 TRANSISTORS), CIRCUIT  
* SIMULATION TIME IS INCREASED.    
*  
* CONNECTIONS:  PLUS  
*                |  ADJUST  
*                |  |  MINUS  
*                |  |  |  
.SUBCKT LM185    1  5  6  
*  
R6 1 2 200E3  
R7 2 3 50E3  
R8 3 4 300E3  
Q14 6 5 4 PNPNOM  
Q13 7 7 1 PNPNOM  
Q10 7 3 8 NPNNOM 10  
Q9 8 12 6 NPNNOM  
Q12 9 7 1 PNPNOM  
Q11 9 2 8 NPNNOM  
R5 1 12 600E3  
Q8 12 12 6 NPNNOM  
Q7 13 9 1 PNPNOM  
Q6 13 12 6 NPNNOM  
R2 1 14 7.5E3  
Q4 15 15 14 PNPNOM  
Q5 15 13 16 NPNNOM  
R3 16 6 500  
Q3 17 15 1 PNPNOM  
R1 17 6 100E3  
Q1 1 17 6 NPNNOM  
C1 17 15 20E-12  
C2 13 9 20E-12  
D1 6 1 DZENER  
.MODEL NPNNOM NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL PNPNOM PNP(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL DZENER D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 6.3
+        IBV = .001
+ )
.ENDS LM185  
*$
*  
* RAD: PRERAD  
* TEMP= -55  
*  
* NOTE: TRR MEASUREMENT WAS MADE @ 10MA/10MA/2.5MA  
*  
*** CAUTION: THE MEASURED TRR AND THE PSPICE CKT. SIMULATED TRR ARE DIFFERENT  
*            THIS COULD POTENTIALLY LEAD TO ERRORS IN CKT. SIMULATIONS IF USED  
*            AS A RECTIFIER OR IN SWITCHING APPLICATIONS.  
*  
* MEASURED TRR = 687.5NS, SIMULATED TRR = 443.1NS.  
*  
*  
.SUBCKT LM185/-55C  99  2  
D1  2   99   DLEAK  
R1  2   99   1E12  
R2  6   99   0.085  
M1  2   2   6   8   MOS1  
R3  6   8   1E12  
D2  99   2   DFOR  
.MODEL DLEAK    D       (
+         IS = 4.5E-6
+         RS = 0.1117427
+          N = 105
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL MOS1     NMOS    (
+      LEVEL = 1
+        VTO = 2.424
+         KP = 1E7
+      GAMMA = 0
+        PHI = .6
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CBD = 0
+        CBS = 0
+         IS = 1E-14
+         PB = .8
+       CGSO = 0
+       CGDO = 0
+       CGBO = 0
+        RSH = 0
+         CJ = 0
+         MJ = .5
+       CJSW = 0
+       MJSW = .33
+         JS = 1E-08
+        TOX = .0000001
+        NSS = 0
+        NFS = 0
+        TPG = 1
+         XJ = 0
+         LD = 0
+         UO = 600
+      UCRIT = 10000
+       UEXP = 0
+       UTRA = 0
+       VMAX = 0
+       NEFF = 1
+        XQC = 1
+         KF = 0
+         AF = 1
+         FC = .5
+      DELTA = 0
+      THETA = 0
+        ETA = 0
+      KAPPA = .2
+ )
.MODEL DFOR     D       (
+         IS = 2.923266E-10
+         RS = 18.800808
+          N = 1.6458985
+         TT = 6.0E-7
+        CJO = 6.732155E-11
+         VJ = 0.6208282
+          M = 0.2203896
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = 0.5
+         BV = 1E5
+        IBV = .001
+ )
.ENDS LM185/-55C
*
*$
*  
* RAD: PRERAD  
* TEMP= 125  
*  
*** NOTE: TRR MEASUREMENT WAS MADE @ 10MA/10MA/2.5MA  
*  
*** CAUTION: THE MEASURED TRR AND THE PSPICE CKT. SIMULATED TRR ARE DIFFERENT  
*            THIS COULD POTENTIALLY LEAD TO ERRORS IN CKT. SIMULATIONS IF USED  
*            AS A RECTIFIER OR IN SWITCHING APPLICATIONS.  
*  
* MEASURED TRR = 1.877US, SIMULATED TRR = 1.233US.  
*  
*  
.SUBCKT LM185/125C  99  2  
D1  2   99   DLEAK  
R1  2   99   1E12  
R2  6   99   0.15  
M1  2   2   6   8   MOS1  
R3  6   8   1E12  
D2  99   2   DFOR  
.MODEL DLEAK    D       (
+         IS = 1E-6
+         RS = 15.831318
+          N = 45
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1E5
+        IBV = .001
+ )
.MODEL MOS1     NMOS    (
+      LEVEL = 1
+        VTO = 2.598
+         KP = 1E4
+      GAMMA = 0
+        PHI = .6
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CBD = 0
+        CBS = 0
+         IS = 1E-14
+         PB = .8
+       CGSO = 0
+       CGDO = 0
+       CGBO = 0
+        RSH = 0
+         CJ = 0
+         MJ = .5
+       CJSW = 0
+       MJSW = .33
+         JS = 1E-08
+        TOX = .0000001
+        NSS = 0
+        NFS = 0
+        TPG = 1
+         XJ = 0
+         LD = 0
+         UO = 600
+      UCRIT = 10000
+       UEXP = 0
+       UTRA = 0
+       VMAX = 0
+       NEFF = 1
+        XQC = 1
+         KF = 0
+         AF = 1
+         FC = .5
+      DELTA = 0
+      THETA = 0
+        ETA = 0
+      KAPPA = .2
+ )
.MODEL DFOR     D       (
+         IS = 1.024781E-8
+         RS = 10.4280679
+          N = 2.1779911
+         TT = 1.6E-6
+        CJO = 7.791736E-11
+         VJ = 0.4
+          M = 0.2944435
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = 0.5
+         BV = 1E5
+        IBV = .001
+ )
.ENDS LM185/125C
*$
* MANUFACTURERS PART NO. = LM185BYH/883  (NATIONAL SEMICONDUCTOR)  
* TYPE: IC_LINEAR  
* SUBTYPE: REFERENCE  
* THIS FILE CONTAINS ONE RADIATION MODEL OF THE 2 TERMINAL 1.2V REF.  
* PARAMETER MODEL EXTRACTED FROM MEASURED DATA  
* CREATION DATE : 07-23-90  
*  
* RAD: 1.13E12  
* TYPE: NEUTRON              
*  
* TEMP= 27  
*  
*** NOTE: TRR MEASUREMENT WAS MADE @ 10MA/10MA/2.5MA  
*  
*** CAUTION: THE MEASURED TRR AND THE PSPICE CKT. SIMULATED TRR ARE DIFFERENT  
*            THIS COULD POTENTIALLY LEAD TO ERRORS IN CKT. SIMULATIONS IF USED  
*            AS A RECTIFIER OR IN SWITCHING APPLICATIONS.  
*  
*  
* MEASURED TRR = 451.250NS, SIMULATED TRR = 360.4NS.  
*  
*  
.SUBCKT LM185/27C/RAD 99  2  
D1  2   99   DLEAK  
R1  2   99   1.001E12  
R2  6   99   0.33  
M1  2   2   6   8   MOS1  
R3  6   8   1E12  
D2  99   2   DFOR  
.MODEL DLEAK    D       (
+         IS = 3E-6
+         RS = 40
+          N = 65
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.MODEL MOS1     NMOS    (
+      LEVEL = 1
+        VTO = 2.558
+         KP = 5E6
+      GAMMA = 0
+        PHI = .6
+     LAMBDA = 0
+         RD = 0
+         RS = 0
+        CBD = 0
+        CBS = 0
+         IS = 1E-14
+         PB = .8
+       CGSO = 0
+       CGDO = 0
+       CGBO = 0
+        RSH = 0
+         CJ = 0
+         MJ = .5
+       CJSW = 0
+       MJSW = .33
+         JS = 1E-08
+        TOX = .0000001
+        NSS = 0
+        NFS = 0
+        TPG = 1
+         XJ = 0
+         LD = 0
+         UO = 600
+      UCRIT = 10000
+       UEXP = 0
+       UTRA = 0
+       VMAX = 0
+       NEFF = 1
+        XQC = 1
+         KF = 0
+         AF = 1
+         FC = .5
+      DELTA = 0
+      THETA = 0
+        ETA = 0
+      KAPPA = .2
+ )
.MODEL DFOR     D       (
+         IS = 6.652648E-9
+         RS = 17.4283533
+          N = 2.0158844
+         TT = 4.8E-7
+        CJO = 6.069386E-11
+         VJ = 0.540285
+          M = 0.2625517
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = 0.4868582
+         BV = 9.9999E+13
+        IBV = .001
+ )
.ENDS LM185/27C/RAD
*$
*
*---------------------------------------------------------------MC7805C
.SUBCKT MC7805C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
* MANUFACTURERS PART NO. = REF02/883/J  (PRECISION MONOLITHIC)
* SUBTYPE: REFERENCE
* THIS FILE CONTAINS 1 PRERAD ROOM TEMPERATURE MACROMODEL OF THE REF02
* PRECISION 5V REFERENCE.
*
*
* PLEASE NOTE THE FOLLOWING:
*
* THIS MODEL IS TO BE USED AT 27 C.
*
*------------------------------------------------------------------------------
*
*
*                IN
*                 |  TEMP
*                 |    |   GND
*                 |    |    |   TRIM
*                 |    |    |    |   OUT
*                 |    |    |    |    |
.SUBCKT REF-02    2   3   4   5   6
R1 11 3 1000
R2 3 4 9353.193
R3 1 7 10000
R4 1 8 10000
R6 1000 2 1000
DR6 1000 1 DR6
.MODEL DR6 D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
RBREF 9 5 .5
Q1 7 9 11 NREF1 8
Q2 8 5 3 NREF1
.MODEL NREF1 NPN (
+         IS = 1E-8
+         BF = 200
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
R7 12 13 100
C1 13 7 .001P
RC1 13 4 100MEG
EA 120 4 8 7 1000
RIN 8 7 100K
RO 12 120 5
ECL 302 4 2 4 1
V+ 301 302 DC 0
DC+ 12 301 DMOD2
VDC 300 4 DC 1
DC- 300 12 DMOD2
.MODEL DMOD2 D (
+         IS = 1E-20
+         RS = 0
+          N = .5
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
RB 200 18 100
DB 200 17 DB
.MODEL DB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
EB 17 4 13 4 1
IBIAS 2 201 .475M
RTEST 200 201 1K
QPASS 16 18 6 NTYPE
.MODEL NTYPE NPN (
+         IS = 1E-16
+         BF = 53.0948
+         NF = 1
+        VAF = 22.6799
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
DPASS 6 16 DMOD
R15 2 16 20
R12 6 5 6.1K
R11 5 4 2K
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.ENDS REF-02
*$
*
*---------------------------------------------------------------UPC7805
.SUBCKT UPC7805 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
*---------------------------------------------------------------SG7805C
.SUBCKT SG7805C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
* MANUFACTURERS PART NO.= SG7805AIG  (SILICON GENERAL)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMP. DEPENDENT MODEL OF THE SG7805
* REGULATOR.
*
*------------------------------------------------------------------------------
*
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT.  IT
* INCLUDES POWER-UP AND POWER-DOWN EFFECTS.
* IT IS NECESSARY TO SET ITL1=300 ITL2=300 WITH THE .OPTIONS COMMAND FOR
* 100%  CONVERGENCE.  THESE SETTINGS DETERMINE THE NUMBER OF ITERATIONS
* ALLOWED FOR  THE CALCULATION OF THE DC AND BIAS PT VALUES WHEN THE
* STARTING POINT IS  CONSIDERED "BLIND" OR AN "EDUCATED GUESS".
* OTHER SETTINGS MAY WORK, BUT HAVE NOT BEEN TESTED YET.
*
*
*
.SUBCKT SG7805  1 2  3
*               |  |   |
*              IN  |   |
*                 OUT  |
*                     GND
*




*** VOLTAGE REFERENCE AND BIAS CURRENT SECTION ***
DZ1  4 1 DZ1
.MODEL DZ1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.5
+        IBV = .001
+ )
RQ   4 17 112090 TC=0.003483, -4.9343E-6
RR   17 18 4.7 TC=0.003449, -5.495E-6
DR   16 18 DR
.MODEL DR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.2651
+        IBV = .001
+ )
RZ 16 18 1MEG
L1 16 3 IND1 0.796M
.MODEL IND1 IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 0.00236
+        TC2 = 1.24436E-5
+ )
*** ERROR AMPLIFIER SECTION ***
EP 22 3 17 15 300
RO 22 6 25
DC- 3 6 DCLAMP
DC+ 6 19 DCLAMP
.MODEL DCLAMP D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
V+ 19 23 DC -1
E+ 23 3 1 3 1
RP 6 7 50
CPZ 7 3 0.5U
*** QUIESCENT CURRENT ***
GB 1 9 17 3 0.5002M
RQUIES 12 3 3396 TC=0.006886, 4.655264E-5
*** SHORT CIRCUIT AND FOLDBACK CURRENT ***
DBL 9 8 DBL
.MODEL DBL D(
+         IS = 1E-4
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
EB 8 3 7 3 2
RC 1 14 0.2
DC 14 13 DC
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1.617
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
RB 9 11 100
QP 13 11 5 QP
.MODEL QP NPN(
+         IS = 1E-12
+         BF = 70K
+         NF = 1
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
DCL 9 10 DCL
.MODEL DCL D(
+         IS = 1E-4
+         RS = 0
+          N = 2
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
QCL 10 20 12 QLIMIT
.MODEL QLIMIT NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
RSC 5 12 0.275 TC=0.001885, 9.363636E-6
RBCL 20 5 1600
RFBCL 1 21 51.17K TC= 0.002528, -1.5164E-5
DZFB 20 21 DZFB
.MODEL DZFB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 15.26
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -9.5474743E-4
+       TBV2 = 1.478994E-5
+       TRS1 = 0
+       TRS2 = 0
+ )
R24 15 3 600
R23 12 15 1800
*** OUTPUT RESISTANCE ***
ROUT 12 2 0.036 TC=0.002616, -1.50463E-5
DDIS 12 1 DMOD
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 0.7
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS SG7805
*$
*
* MANUFACTURERS PART NO.= SG7805AIG  (SILICON GENERAL)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD 27 C TEMPERATURE MACROMODEL
* OF THE SG7805AIG REGULATOR.
*
*---------------------------------------------------------------------------
* PLEASE NOTE THE FOLLOWING:
*
* 1) THIS MODEL IS TO BE USED FOR ROOM TEMPERATURE SIMULATIONS.  THE
*  SPICE TEMPERATURE CORRECTIONS WILL NOT WORK.
*
*
*
.SUBCKT SG7805/27C  1  2   3
*                   |  |   |
*                  IN  |   |
*                     OUT  |
*                        GND
DZ1 16 1 DZ1
.MODEL DZ1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 0.75
+        IBV = .001
+ )
RQ 16 17 113K
RR 17 18 7.0476
DR 3 18 DR
.MODEL DR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.27
+        IBV = .001
+ )
RDR 3 17 30K
GQ 1 4 17 3 1M
ER 4 3 17 3 1
RIN 4 15 100MEG
RC 1 14 0.2
DBK 14 13 DBK
.MODEL DBK D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
EP 19 3 4 15 250
RO 19 6 25
DC- 3 6 DC
DC 6 20 DC
.MODEL DC D(
+         IS = 1E-20
+         RS = 0
+          N = 0.1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
EC 20 3 1 3 1
RP 6 7 75
RPZ 7 8 0.1
CPZ 8 3 0.1U
GB 1 9 17 3 2.184M
EB 22 3 7 3 1
DB1 9 22 DB1
.MODEL DB1 D(
+         IS = 1E-14
+         RS = 0
+          N = 0.01
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
CDB1 9 22 10U
RB1 9 10 1
RB2 10 11 750
RBC 12 11 7500
CBC 13 12 0.002U
CBE 11 21 0.001U
QP 13 11 5 QP
.MODEL QP NPN(
+         IS = 1E-16
+         BF = 2296
+         NF = 1
+        VAF = 50
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
QLIMIT 10 23 21 QLIMIT
.MODEL QLIMIT NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
RBC1 23 5 2400
RSENSE 5 21 0.2303
RFBL 1 24 80K
DZFB 23 24 DZFB
.MODEL DZFB D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 14.07
+        IBV = .001
+ )
RFB1 15 3 6K
RFB2 21 15 18K
ROUT 21 2 0.04
.ENDS SG7805/27C
*$
*
*---------------------------------------------------------------UC7805C
.SUBCKT UC7805C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
*---------------------------------------------------------------LM7812C
.SUBCKT LM7812C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------uA7812C
.SUBCKT UA7812C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------LAS1512
.SUBCKT LAS1512 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------MC7812C
.SUBCKT MC7812C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------UPC7812
.SUBCKT UPC7812 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------SG7812C
.SUBCKT SG7812C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
* MANUFACTURERS PART NO.= SG7812AIG  (SILICON GENERAL)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMP. DEPENDENT MODEL OF THE SG7812
* REGULATOR
*
*------------------------------------------------------------------------------
*
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT.  IT
* INCLUDES POWER-UP AND POWER-DOWN EFFECTS.
* IT IS NECESSARY TO SET ITL1=300 ITL2=300 WITH THE .OPTIONS COMMAND FOR
* 100%  CONVERGENCE.  THESE SETTINGS DETERMINE THE NUMBER OF ITERATIONS
* ALLOWED FOR  THE CALCULATION OF THE DC AND BIAS PT VALUES WHEN THE
* STARTING POINT IS  CONSIDERED "BLIND" OR AN "EDUCATED GUESS".
* OTHER SETTINGS MAY WORK, BUT HAVE NOT BEEN TESTED YET.
*
*
*
.SUBCKT SG7812  1 2  3
*               |  |   |
*              IN  |   |
*                 OUT  |
*                     GND
*
*** VOLTAGE REFERENCE AND BIAS CURRENT SECTION ***
DZ1  4 1 DZ1
.MODEL DZ1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 0.75
+        IBV = .001
+ )
RQ   4 17 86343.84 TC=5.3597E-4, 5.0408E-5
RR   17 18 5.2447 TC=0.005772, 6.2073E-5
DZR   16 18 DR
.MODEL DR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.2588
+        IBV = .001
+ )
RZ 16 18 1MEG
L1 16 3 IND1 0.3573M
.MODEL IND1 IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 0.001123
+        TC2 = 6.8566E-5
+ )
*** ERROR AMPLIFIER SECTION ***
EA 22 3 17 15 300
ROUT 22 6 10
D- 3 6 DCLAMP
D+ 6 19 DCLAMP
.MODEL DCLAMP D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
V+ 19 23 DC -1
E+ 23 3 1 3 1
RP 6 7 500
CP 7 3 CAP1 0.1U
.MODEL CAP1 CAP(
+          C = 1
+        VC1 = 0
+        VC2 = 0
+        TC1 = -0.002
+        TC2 = 1E-4
+ )
*** QUIESCENT CURRENT ***
GB 1 9 17 3 0.4944M
RQUIES 12 3 10572.61 TC=0.013985, 1.28953E-4
*** SHORT CIRCUIT AND FOLDBACK CURRENT ***
DBL 9 8 DBL
.MODEL DBL D(
+         IS = 1E-4
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
EB 8 3 7 3 2
RC 1 14 0.2
DC 14 13 DC
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1.6339
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
RB 9 11 100
QP 13 11 5 QP
.MODEL QP NPN(
+         IS = 1E-12
+         BF = 70K
+         NF = 1
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
DCL 9 10 DCL
.MODEL DCL D(
+         IS = 1E-4
+         RS = 0
+          N = 2
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
QCL 10 20 12 QCL
.MODEL QCL NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
RSC 5 12 0.578 TC=0.00131, 1.2433E-5
RBCL 20 5 200
RFB 1 21 6.17043K TC=0.001143, -1.081421E-5
DZFB 20 21 DZFB
.MODEL DZFB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 14.79
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -1.78236E-4
+       TBV2 = 4.2164E-6
+       TRS1 = 0
+       TRS2 = 0
+ )
R24 15 3 600
R23 12 15 5160
*** OUTPUT RESISTANCE ***
RO 12 2 0.02 TC=-8.3333E-4, -4.1667E-5
DDIS 2 1 DMOD
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 0.7
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS SG7812
*$
*
* MANUFACTURERS PART NO.= SG7812AIG  (SILICON GENERAL)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD 27 C TEMPERATURE  MODEL
* OF THE SG7812 REGULATOR.
*
*
*---------------------------------------------------------------------------
* PLEASE NOTE THE FOLLOWING:
*
*
* 1) THIS MODEL IS TO BE USED FOR ROOM TEMPERATURE SIMULATIONS.  THE
*    SPICE TEMPERATURE CORRECTIONS WILL NOT WORK.
*
*
*----------------------------------------------------------------
*
*
.SUBCKT SG7812/27C  1  2   3
*                   |  |   |
*                  IN  |   |
*                     OUT  |
*                        GND
*
DZ1 16 1 DZ1
.MODEL DZ1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 0.75
+        IBV = .001
+ )
RQ 16 17 113K
RR 17 18 7.0476
DR 3 18 DR
.MODEL DR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.27
+        IBV = .001
+ )
RDR 3 17 30K
GQ 1 4 17 3 1M
ER 4 3 17 3 1
RIN 4 15 100MEG
RC 1 14 0.2
DBK 14 13 DBK
.MODEL DBK D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
EP 19 3 4 15 250
RO 19 6 25
DC- 3 6 DC
DC 6 20 DC
.MODEL DC D(
+         IS = 1E-20
+         RS = 0
+          N = 0.1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
EC 20 3 1 3 1
RP 6 7 75
RPZ 7 8 0.1
CPZ 8 3 0.1U
GB 1 9 17 3 2.184M
EB 22 3 7 3 1
DB1 9 22 DB1
.MODEL DB1 D(
+         IS = 1E-14
+         RS = 0
+          N = 0.01
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
CDB1 9 22 10U
RB1 9 10 1
RB2 10 11 750
RBC 12 11 7500
CBC 13 12 0.002U
CBE 11 21 0.001U
QP 13 11 5 QP
.MODEL QP NPN(
+         IS = 1E-16
+         BF = 2296
+         NF = 1
+        VAF = 50
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
QLIMIT 10 23 21 QLIMIT
.MODEL QLIMIT NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
RBC1 23 5 2400
RSENSE 5 21 0.7285
RFBL 1 24 57.6K
DZFB 23 24 DZFB
.MODEL DZFB D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 14.07
+        IBV = .001
+ )
RFB1 15 3 6K
RFB2 21 15 51.6K
ROUT 21 2 1E-6
.ENDS SG7812/27C
*$
*
*---------------------------------------------------------------UC7812C
.SUBCKT UC7812C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------LM7815C
.SUBCKT LM7815C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
*---------------------------------------------------------------uA7815C
.SUBCKT UA7815C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
* MANUFACTURERS PART NO. = UA78M05HM   (FAIRCHILD)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD MODEL AT 27 C OF THE LM7805 THAT WAS
* DEVELOPED  UNDER THE GUIDANCE OF GREGORY M. WIERZBA AT MICHIGAN STATE
* UNIVERSITY
*
* PLEASE NOTE THE FOLLOWING:
*
*   1) THIS MODEL IS TO BE USED FOR ROOM TEMPERATURE SIMULATIONS. THE BUILT-
*      IN  SPICE TEMPERATURE CORRECTIONS WILL NOT WORK.
*   2) RIPPLE REJECTION, OUTPUT IMPEDANCE, LINE TRANSIENT, AND LOAD
*      TRANSIENT RESPONSE ARE MODELED BASED ON LABORATORY
*      MEASUREMENTS.  THE CORRELATION IS QUITE GOOD. THE SIMULATION VALUES
*      ARE WITHIN THE PRODUCT SPEC LIMITS.
*   3) CURRENT LIMITING IS CURRENTLY SET FOR 600MA WITH FOLDBACK EFFECTS
*      FOR  SAFE OPERATING REGION, BUT IF THIS CAUSES PROBLEMS IT CAN EASILY
*      BE  CHANGED TO A HIGHER LEVEL FOR THE USER.
*   4) QUIESCENT CURRENT HAS ALSO BEEN MODELED BUT REQUIRES MORE LAB
*      VERIFICATION.  DROPOUT AND POWER UP CHARACTERISTICS HAVE NOT BEEN
*      DEVELOPED YET IN THIS MODEL.
*   5) FOR FURTHER DETAILS AND THE MODEL DERIVATION, OBTAIN A COPY OF
*      "CA3085,  LM7805, LM7812, LM7905, LM137 MACROMODEL DEVELOPMENT" BY G. M.
*      WIERZBA  DATED 3/25/91.
*
*
*
*
.SUBCKT UA78M05  1   2    3        99
*               IN   |    |         |
*                   OUT   |         |
*                        GND(PIN)   |
*                               ZERO REFERENCE(EXTERNAL GND)
IBIAS   1 4 3M
VREF    15 3 DC 3.7
ELREG   4 15 1 3 .074M
RIN     4 5 10000
RC      1 14 0.2
EP      6 3 4 5 1200
RP      6 7 10000
RZ      7 8 10
CPZ     8 3 10U
EB      16 3 7 3 1
DLIM    9 16 DMOD
CBYPASS 9 16 100U
RB      9 11 26
RBC     12 11 400
CBC     13 12 0.001U
QPASS   13 11 2 QMOD
DBK     14 13 DMOD
RFB1    2 5 1756.5
RFB2    5 3 5000
GLIMIT  3 9 POLY(1) 13 2 .6279M -5.5186U
GFB     9 3 POLY(1) 18 99 0 15.1775U
EFB     17 99 1 2 1
DZFB    18 17 DZ
.MODEL DZ D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.5
+        IBV = .001
+ )
RFB     18 99 1K
.MODEL QMOD NPN (
+         IS = 1E-16
+         BF = 1000
+         NF = 1
+        VAF = 100
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL DMOD D (
+         IS = 30F
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.ENDS UA78M05
*$
*
* MANUFACTURERS PART NO. = UA78M12HM   (FAIRCHILD)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD MODEL AT 27 C OF THE LM7812 THAT WAS
* DEVELOPED UNDER THE GUIDANCE OF GREGORY M. WIERZBA AT
* MICHIGAN STATE UNIVERSITY.
*
* PLEASE NOTE THE FOLLOWING:
*   1) THIS MODEL IS TO BE USED FOR ROOM TEMPERATURE SIMULATIONS. THE BUILT-
*      IN  SPICE TEMPERATURE CORRECTIONS WILL NOT WORK.
*   2) RIPPLE REJECTION, OUTPUT IMPEDANCE, LINE TRANSIENT, AND LOAD
*      TRANSIENT  RESPONSE ARE MODELED BASED ON LABORATORY
*      MEASUREMENTS.  THE CORRELATION  IS QUITE GOOD. THE SIMULATION VALUES
*      ARE WITHIN THE PRODUCT SPEC LIMITS.
*   3) CURRENT LIMITING IS CURRENTLY SET FOR 600MA WITH FOLDBACK EFFECTS
*      FOR  SAFE OPERATING REGION, BUT IF THIS CAUSES PROBLEMS IT CAN EASILY
*      BE  CHANGED TO A HIGHER LEVEL FOR THE USER.
*   4) QUIESCENT CURRENT HAS ALSO BEEN MODELED BUT REQUIRES MORE LAB
*      VERIFICATION.  DROPOUT AND POWER UP CHARACTERISTICS HAVE NOT BEEN
*      DEVELOPED YET IN THIS MODEL.
*   5) FOR FURTHER DETAILS AND THE MODEL DERIVATION, OBTAIN A COPY OF
*      "CA3085,  LM7805, LM7812, LM7905, LM137 MACROMODEL DEVELOPMENT" BY G. M.
*      WIERZBA  DATED 3/25/91.
*
.SUBCKT UA78M12/27C  1   2   3       99
*                   IN   |   |       |
*                       OUT  |       |
*                           GND(PIN) |
*                                   ZERO REFERENCE(EXTERNAL GND)
IBIAS   1 4 3M
VREF    15 3 DC 3.7
ELREG   4 15 1 3 0.3083M
RIN     4 5 10000
RC      1 14 0.2
EP      6 3 4 5 1200
RP      6 7 10000
RZ      7 8 10
CPZ     8 3 0.01U
EB      16 3 7 3 1
DLIM    9 16 DMOD
CBYPASS 9 16 100U
RB      9 11 26
RBC     12 11 400
CBC     13 12 0.001U
QPASS   13 11 2 QMOD
DBK     14 13 DMOD
RFB1    2 5 11216.2162
RFB2    5 3 5000
GLIMIT  3 9 POLY(1) 13 2 .6279M -5.5186U
GFLDBCK 9 3 POLY(1) 18 99 0 14U
EFB     17 99 13 2 1
DFB     18 17 DZ
.MODEL DZ D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.5
+        IBV = .001
+ )
RFB     18 99 1K
.MODEL QMOD NPN (
+         IS = 1E-16
+         BF = 1000
+         NF = 1
+        VAF = 100
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL DMOD D (
+         IS = 30F
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.ENDS UA78M12/27C
*$
*
* MANUFACTURERS PART NO. = UA78M15HM   (FAIRCHILD)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMP. DEPENDENT MODEL OF THE UA78M15
* REGULATOR
*
*------------------------------------------------------------------------------
*
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT.  IT
* INCLUDES POWER-UP AND POWER-DOWN EFFECTS.
* IF IT IS NECESSARY, SET ITL1=300 ITL2=300 WITH THE .OPTIONS COMMAND FOR
* 100%  CONVERGENCE.  THESE SETTINGS DETERMINE THE NUMBER OF ITERATIONS
* ALLOWED FOR  THE CALCULATION OF THE DC AND BIAS PT VALUES WHEN THE
* STARTING POINT IS  CONSIDERED "BLIND" OR AN "EDUCATED GUESS".
* OTHER SETTINGS MAY WORK, BUT HAVE NOT BEEN TESTED YET.
*
*
*
.SUBCKT UA78M15  1  2   3
*                |  |   |
*               IN  |   |
*                  OUT  |
*                      GND
*
*** VOLTAGE REFERENCE AND BIAS CURRENT SECTION ***
DZ1  4 1 DZ1
.MODEL DZ1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 0.75
+        IBV = .001
+ )
RQ   4 17 86343.84 TC=5.3597E-4, 5.0408E-5
RR   17 18 5.2447 TC=0.005772, 6.2073E-5
DZR   16 18 DR
.MODEL DR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.2588
+        IBV = .001
+ )
RZ 16 18 1MEG
L1 16 3 IND1 .3573M
.MODEL IND1 IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 0.001123
+        TC2 = 6.8566E-5
+ )
*** ERROR AMPLIFIER SECTION ***
EA 22 3 17 15 300
ROUT 22 6 10
D- 3 6 DCLAMP
D+ 6 19 DCLAMP
.MODEL DCLAMP D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
V+ 19 23 DC -1
E+ 23 3 1 3 1
RP 6 7 500
CP 7 3 CAP1 0.1U
.MODEL CAP1 CAP(
+          C = 1
+        VC1 = 0
+        VC2 = 0
+        TC1 = -0.002
+        TC2 = 1E-4
+ )
*** QUIESCENT CURRENT ***
GB 1 9 17 3 0.4944M
RQUIES 12 3 7213 TC=0.013985, 1.28953E-4
*** SHORT CIRCUIT AND FOLDBACK CURRENT ***
DBL 9 8 DBL
.MODEL DBL D(
+         IS = 1E-4
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
EB 8 3 7 3 2
RC 1 14 0.2
DC 14 13 DC
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1.6339
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
RB 9 11 100
QP 13 11 5 QP
.MODEL QP NPN(
+         IS = 1E-12
+         BF = 70K
+         NF = 1
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
DCL 9 10 DCL
.MODEL DCL D(
+         IS = 1E-4
+         RS = 0
+          N = 2
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
QCL 10 20 12 QCL
.MODEL QCL NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
RSC 5 12 1.2721 TC=0.00131, 1.2433E-5
RBCL 20 5 200
RFB 1 21 6089 TC=0.001143, -1.081421E-5
DZFB 20 21 DZFB
.MODEL DZFB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 10
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -1.78236E-4
+       TBV2 = 4.2164E-6
+       TRS1 = 0
+       TRS2 = 0
+ )
R24 15 3 600
R23 12 15 6900
*** OUTPUT RESISTANCE ***
RO 12 2 0.02 TC=-8.3333E-4, -4.1667E-5
DDIS 2 1 DMOD
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 0.7
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS UA78M15
*$
*
* MANUFACTURERS PART NO. = UA79M05HM   (FAIRCHILD)
* SUBTYPE: REGULATOR
*
* THIS FILE CONTAINS A PRE-RAD MODEL AT 27 C OF THE LM7905 THAT WAS
* DEVELOPED UNDER THE GUIDANCE OF GREGORY M. WIERZBA AT
* MICHIGAN STATE UNIVERSITY.

* PLEASE NOTE THE FOLLOWING:
*   1) THIS MODEL IS TO BE USED FOR ROOM TEMPERATURE SIMULATIONS. THE BUILT-
*       IN  SPICE TEMPERATURE CORRECTIONS WILL NOT WORK.
*   2) RIPPLE REJECTION, OUTPUT IMPEDANCE, LINE TRANSIENT, AND LOAD
*       TRANSIENT  RESPONSE ARE MODELED BASED ON LABORATORY
*       MEASUREMENTS.  THE CORRELATION  IS QUITE GOOD. THE SIMULATION VALUES
*       ARE WITHIN THE PRODUCT SPEC LIMITS.
*   3) CURRENT LIMITING IS CURRENTLY SET FOR 600MA WITH FOLDBACK EFFECTS
*       FOR  SAFE OPERATING REGION, BUT IF THIS CAUSES PROBLEMS IT CAN EASILY
*       BE  CHANGED TO A HIGHER LEVEL FOR THE USER.
*   4) QUIESCENT CURRENT HAS ALSO BEEN MODELED BUT REQUIRES MORE LAB
*      VERIFICATION.  DROPOUT AND POWER UP CHARACTERISTICS HAVE NOT BEEN
*      DEVELOPED YET IN THIS MODEL.
*   5) FOR FURTHER DETAILS AND THE MODEL DERIVATION, OBTAIN A COPY OF
*      "CA3085,  LM7805, LM7812, LM7905, LM137 MACROMODEL DEVELOPMENT" BY G. M.
*       WIERZBA  DATED 3/25/91.
*
*
*
*
.SUBCKT UA79M05  1        2     3     99
*               GND(PIN)  |     |     |
*                        OUT    |     |
*                              IN     |
*                                ZERO REFERENCE(EXTERNAL GND)
VREF    1 11 DC 3.7
ELREG   11 4 1 3 0.00234
IBIAS   4 3 DC 3.5M
RIN     4 5 10000
E1      6 3 5 4 1000
RP      6 7 50000
C1      7 3 0.01U
E2      12 3 7 3 1
DLIMIT  9 12 DMOD
GLIMIT  3 9 POLY (1) 2 3 0.4M -4.3U
GFB     9 3 POLY (1) 16 99 -0.2M 0.015M
EFB     15 99 2 3 1
DFB     16 15 DZ
RFB     16 99 1000
R1      5 10 1.7568K
R2      1 5 5K
RB      9 8 5
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.MODEL DZ D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.5
+        IBV = .001
+ )
QOUT    10 8 3 QMOD
.MODEL QMOD NPN (
+         IS = 1E-14
+         BF = 1000
+         NF = 1
+        VAF = 100
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
RCQ     10 14 1000
CQ     14 8 0.0001U
RZOUT    10 2 0.04
.ENDS UA79M05
*$
*
* MANUFACTURERS PART NO. = UA79M15HM   (FAIRCHILD)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMP. DEPENDENT MODEL OF THE UA79M15
* REGULATOR
*
*------------------------------------------------------------------------------
*
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT.  IT
* INCLUDES POWER-UP AND POWER-DOWN EFFECTS.   IT IS NECESSARY TO SET
* ITL1=300 ITL2=300 WITH THE  .OPTIONS COMMAND FOR 100% CONVERGENCE.
* THESE SETTINGS DETERMINE THE  NUMBER OF ITERATIONS ALLOWED FOR THE
* CALCULATION OF THE DC AND BIAS PT  VALUES WHEN THE STARTING POINT IS
* CONSIDERED "BLIND" OR AN "EDUCATED GUESS".  OTHER SETTINGS MAY WORK,
* BUT HAVE NOT BEEN TESTED YET.
*
*
.SUBCKT UA79M15  1       2   3   99
*                |       |   |    |
*              GND(PIN)  |   |    |
*                       OUT  |    |
*                           IN  ZERO REFERENCE(EXTERNAL GND)
*
*** VOLTAGE REFERENCE SECTION ***
LZR 4 1 IND1 0.2079M
.MODEL IND1 IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 0.021188
+        TC2 = 3.9548E-4
+ )
DZR  29 4 DZR
.MODEL DZR D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 2.7117
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -2.4708E-5
+       TBV2 = 3.1346E-7
+       TRS1 = 0
+       TRS2 = 0
+ )
RZR 29 4 1MEG
RR   29 15 5.8475 TC=0.013783, 2.0804E-4
RQ   15 22 42072.4191 TC=0.007522, 1.3907E-4
D1   3 22 D1
.MODEL D1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 2
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -0.004583
+       TBV2 = 2.08333E-5
+       TRS1 = 0
+       TRS2 = 0
+ )
****
FQ 1 3 POLY(3) VQ1 VQ2 VQ3 0 1 1 -1
*** ERROR AMPLIFIER SECTION ***
EA 9 3 5 15 600
RO 6 9 200
D+ 6 20 DC
E+ 20 21 1 3 1
V+ 21 3 -1
D- 19 6 DC
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
V- 19 3 DC 1
***
RP 6 7 1
CP 7 3 1U
*** QUIESCENT CURRENT SECTION ***
EQ1 23 99 TABLE {V(1,3)} (2,0) (6.5,4.5)
VQ1 23 24 DC 0
RQ1 24 99 2251.1256 TC=0.004046, 1.1071E-5
EQ2 25 99 TABLE {V(1,3)} (6.5,0) (16,9.5)
VQ2 25 26 DC 0
RQ2 26 99 5757.81 TC=0.008862, 5.369E-5
EQ3 27 99 TABLE {V(1,3)} (16,0) (16.5,0.5)
VQ3 27 28 DC 0
RQ3 289 155.4 TC=0.005318, 1.2798E-5
***
GB 1 8 1 15 4M
GCOMP 3 1 1 15 4M
DB 8 18 DB
.MODEL DB D(
+         IS = 1E-14
+         RS = 0.1
+          N = 0.1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
EB 18 3 7 3 1
RB 8 10 10
*** CURRENT LIMIT AND FOLDBACK CURRENT SECTION ***
QL 1 14 14 QTEMP
.MODEL QTEMP NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
RFB 12 14 34.829K TC=0.003476, -3.2976E-6
DZFB 13 12 DZFB
.MODEL DZFB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 7.8523
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -0.001336
+       TBV2 = 9.3921E-6
+       TRS1 = 0
+       TRS2 = 0
+ )
QCL 10 13 3 QMOD
RBCL 13 17 1K
RCL 17 3 1.19625 TC=6.659E-4, 7.318E-6
***
RBC  11 14 351
CBC  10 11 1N
*** OUTPUT TRANSISTOR ***
QP 16 10 17 QMOD
.MODEL QMOD NPN(
+         IS = 1E-14
+         BF = 70000
+         NF = 1
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
DDO  14 30 DDO
.MODEL DDO D(
+         IS = 1E-14
+         RS = 0
+          N = 1.0876
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
RDDO 30 16 0.1
R23 1 5 2.69K
R22 5 14 12.5K
ROUT 14 2 0.4 TC=0.003976, -2.8869E-5
DDIS 3 14 DDIS
.MODEL DDIS D(
+         IS = 1E-12
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS UA79M15
*$
*
*---------------------------------------------------------------LAS1515
.SUBCKT LAS1515 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
*---------------------------------------------------------------MC7815C
.SUBCKT MC7815C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
*---------------------------------------------------------------SG7815C
.SUBCKT SG7815C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
*---------------------------------------------------------------UC7815C
.SUBCKT UC7815C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
*---------------------------------------------------------------LM140-5
.SUBCKT LM140-5 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
*---------------------------------------------------------------LM140-12
.SUBCKT LM140-12 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------LM140-15
.SUBCKT LM140-15 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
*---------------------------------------------------------------LM140A-5
.SUBCKT LM140A-5 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
*---------------------------------------------------------------LM140A-12
.SUBCKT LM140A-12 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------LM140A-15
.SUBCKT LM140A-15 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
*---------------------------------------------------------------LM340-5
.SUBCKT LM340-5 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
*---------------------------------------------------------------SG340-5
.SUBCKT SG340-5 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
*---------------------------------------------------------------LM340-12
.SUBCKT LM340-12 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------SG340-12
.SUBCKT SG340-12 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------LM340-15
.SUBCKT LM340-15 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
*---------------------------------------------------------------LM340A-5
.SUBCKT LM340A-5 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
*---------------------------------------------------------------TL780-05C
.SUBCKT TL780-05C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=1665, R1_Value=1020
.ENDS
*$
*
*---------------------------------------------------------------LM340A-12
.SUBCKT LM340A-12 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------TL780-12C
.SUBCKT TL780-12C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=694, R1_Value=2448
.ENDS
*$
*
*---------------------------------------------------------------LM340A-15
.SUBCKT LM340A-15 Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*
*---------------------------------------------------------------TL780-15C
.SUBCKT TL780-15C Input Output Ground
   x1 Input Output Ground x_LM78XX PARAMS:
+     Av_feedback=550, R1_Value=3060
.ENDS
*$
*------------------------------------------------------------------------

*** Voltage regulators (positive/adjustable)
*
* LM117 voltage regulator "macromodel" subcircuit
* created using Parts release 5.3 on 04/08/93 at 11:33
* PARTS is a MicroSim product.
*
* connections:     input
*                  |  adjustment pin
*                  |  |   output
*                  |  |   |
.SUBCKT LM117     IN ADJ OUT
*
* POSITIVE ADJUSTABLE VOLTAGE REGULATOR
*
JADJ IN ADJ ADJ JADJMOD ;ADJUSTMENT PIN CURRENT
VREF 4 ADJ 1.25
DBK IN 13 DMOD
*
* ZERO OF RIPPLE REJECTION
*
CBC 13 15 8e-010
RBC 15 5 1000
*
QPASS 13 5 OUT QPASSMOD
RB1 7 6 1
RB2 6 5 128.3
*
* CURRENT LIMITING
*
DSC 6 11 DMOD
ESC 11 OUT VALUE {5.646-0.1125*V(6,5)*V(13,5)}
*
* FOLDBACK CURRENT
*
DFB 6 12 DMOD
EFB 12 OUT VALUE {7.886-0.3727*V(13,5)+0.005097*V(13,5)*V(13,5)
+ -0.02*V(13,5)*V(6,5)}
*
EB 7 OUT 8 OUT 7.691
*
* ZERO OF OUTPUT IMPEDANCE
*
RP 9 8 100
CPZ 10 OUT 3.979e-006
*
DPU 10 OUT DMOD ;POWER-UP CLAMPLING DIODE
RZ 8 10 0.1
EP 9 OUT 4 OUT 100
RI OUT 4 100MEG
*
.MODEL QPASSMOD NPN (IS=30F BF=50 VAF=8.891 NF=2.612)
.MODEL JADJMOD NJF (BETA=5e-005 VTO=-1)
.MODEL DMOD D (IS=30F N=2.612)
.ENDS
*$
*
* MANUFACTURERS PART NO.= LM117HVH  (NATIONAL SEMICONDUCTOR)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT MODEL OF THE
* LM117HVH  THAT WAS DEVELOPED BY GREGORY M. WIERZBA OF MICHIGAN STATE
* UNIVERSITY
*
* PLEASE NOTE THE FOLLOWING:
*
*   1) THIS MODEL CAN BE USED WITH THE .TEMP STATEMENT FOR TEMPERATURE
*      SIMULATIONS.
*   2) THE RIPPLE REJECTION AND LINE TRANSIENT RESPONSE DATA FOUND IN THE
*      NATIONAL DATA SHEET ARE REPORTED BY THE MODEL DEVELOPER TO BE
*      INCORRECT.
*   3) THIS MODEL SIMULATES SLOW POWER-UP TRANSIENTS( RISE TIME > 5US )
*       QUITE   WELL.  A THERMAL OVERLOAD PROTECTOR SHUTS OFF THE REGULATOR
*       DUE TO A  FAST RISING INPUT WITH A DELAY OF APPROXIMATELY 150USEC.
*       THIS IS NOT SIMULATED IN THE MODEL.
*   4) FOR FURTHER DETAILS AND THE MODEL DERIVATION, OBTAIN A COPY OF
*       LM117HVH MACROMODEL DEVELOPMENT" BY G. M. WIERZBA DATED 10/25/90.
*
*** PLEASE NOTE: THE LM117 IS A 1.2 V TO 37 V DEVICE, WHEREAS THE LM117HVH
*                IS A 1.2 V TO 57 V DEVICE. CHANGE THE NECESSARY PARAMETERS
*                BEFORE USING THIS MODEL FOR THE LM117
*
**** PLEASE NOTE THE FOLLOWING 'WORK AROUND' IF OSCILLATIONS OCCUR WITH A
*    CAPACITOR ON THE OUTPUT:
*
*  SERIES VOLTAGE REGULATORS CONTAIN HIGH GAIN FEEDBACK AMPLIFIERS.  AS
*  WITH ANY FEEDBACK CIRCUIT, DRIVING CAPACITIVE LOADS CAN CAUSE
*  INSTABILITY.
*  THE DATA SHEET FOR THE LM117HVH POINTS OUT THAT EVEN 500 PF CAN CAUSE
*  OSCILLATIONS.  ADDING MORE CAPACITANCE, IN GENERAL, MAKES THE PROBLEM
*  WORSE.  THE DATA SHEET SUGGESTS ADDING A LARGE VALUED ELECTROLYTIC OR
*  TANTALUM CAPACITOR TO SUPPRESS THE OSCILLATIONS.  THIS WORKS BECAUSE
*  THE  EFFECTIVE SERIES RESISTANCE (ESR) OF THESE CAPACITORS IS HIGH AND
*  PRODUCES POLE-ZERO CANCELLATION MUCH LIKE THE SERIES RC CIRCUIT
*  ACROSS  A HIGH PERFORMANCE OPAMP INPUT.
*
*  THE FORMULA FOR ESR IN OHMS IS ESR=(DISSIPATION FACTOR)/(2*PI*F*C). SINCE
*  THE DISSIPATION FACTOR IS FAIRLY CONSTANT, THIS RESISTOR IS A NONLINEAR
*  FUNCTION OF FREQUENCY.  THIS IS DIFFICULT TO MODEL IN SPICE.  HOWEVER,
*  MODELING THE CAPACITOR ACCURATELY AT 40 KHZ IS CRITICAL FOR STABILITY BE-
*  CAUSE OF THE EXISTENCE OF A POLE IN THE RIPPLE REJECTION AT THIS
*  FREQUENCY
*
*  THE LM117 MODEL IS STABLE WITH CAPACITIVE LOADS PROVIDED THAT THE ESR IS
*  INCLUDED.  FOR EXAMPLE, IF A 1 OHM RESISTOR IS ADDED IN SERIES WITH A 1 UF
*  LOAD THEN THE TRANSIENTS DIE OUT WITH TIME.  IF THE LOAD CAPACITANCE IS
*  0.1 UF THEN R SHOULD BE 10 OHMS IN ORDER TO MAINTAIN THE SAME DISSIPATION
*  FACTOR.
*
*
*
.SUBCKT LM117HV  1   2   3   111


*                |   |   |    |
*                IN  |   |    |
*                   OUT  |    |
*                       ADJ   |
*                            GND(REFERENCE)
GADJ 1 4 POLY(1) 100 111 48.4U 1.05739E-7 -5.3237E-10
EREF 4 3 POLY(1) 100 111 1.2782 -6.95011E-7 -1.26005E-6 -6.1947E-9
RC 1 14 0.742
DBK 14 13 DLM117HV
CBC 13 15 2.479N
CPZ 10 2 0.796U
HRBC 15 202 POLY(2) VRBC VTJ 0 247 0 0 1.3722
VRBC 202 5 DC 0
QP 13 5 2 QLM117HV
HRB2 5 203 POLY(2) VRB2 VTJ 0 124 0 0 0.68888
VRB2 203 6 DC 0
DSC 6 11 DLM117HV
ESC 11 2 POLY(2) (13,5) (6,5) 2.85 0 0 0 -70.1M
DFB 6 12 DLM117HV
EFB 12 2 POLY(2) (13,5) (6,5) 3.92 -135M 0 1.21M -70.1M
RB1 7 6 1
EB 7 2 8 2 2.56
RZ 8 10 .104
RP 9 8 100
EP 9 2 4 2 103.6
RI 2 4 100MEG
.MODEL QLM117HV NPN (
+         IS = 30F
+         BF = 50
+         NF = 1.604
+        VAF = 14.97
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL DLM117HV D (
+         IS = 30F
+         RS = 0
+          N = 1.604
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
******THERMAL SENSING CIRCUITRY**************
GPD 102 100 POLY(2) (1,2) (1,14) 0 0 0 0 1.347709
RJC 100 101 12
RCA 101 102 12.5
CJA 100 102 0.001
EAMB 102 111 103 111 1
IAMB 111 103 DC 1
RT1 103 104 100 TC=0.01
RT2 104 111 -100.0000001
ETJ 105 111 100 0 1
VTJ 105 106 DC 0
RTJ 106 111 1
.ENDS LM117HV
*$
* LM138 voltage regulator "macromodel" subcircuit
* created using Parts release 5.3 on 04/08/93 at 11:59
* PARTS is a MicroSim product.
*
* connections:     input
*                  |  adjustment pin
*                  |  |   output
*                  |  |   |
.SUBCKT LM138     IN ADJ OUT
*
* POSITIVE ADJUSTABLE VOLTAGE REGULATOR
*
JADJ IN ADJ ADJ JADJMOD ;ADJUSTMENT PIN CURRENT
VREF 4 ADJ 1.24
DBK IN 13 DMOD
*
* ZERO OF RIPPLE REJECTION
*
CBC 13 15 8e-010
RBC 15 5 1000
*
QPASS 13 5 OUT QPASSMOD
RB1 7 6 1
RB2 6 5 128.3
*
* CURRENT LIMITING
*
DSC 6 11 DMOD
ESC 11 OUT VALUE {20.53-0.5*V(6,5)*V(13,5)}
*
* FOLDBACK CURRENT
*
DFB 6 12 DMOD
EFB 12 OUT VALUE {30.11-1.803*V(13,5)+0.02919*V(13,5)*V(13,5)
+ -0.5*V(13,5)*V(6,5)}
*
EB 7 OUT 8 OUT 22.37
*
* ZERO OF OUTPUT IMPEDANCE
*
RP 9 8 100
CPZ 10 OUT 1.326e-005
*
DPU 10 OUT DMOD ;POWER-UP CLAMPLING DIODE
RZ 8 10 0.1
EP 9 OUT 4 OUT 100
RI OUT 4 100MEG
*
.MODEL QPASSMOD NPN (IS=30F BF=50 VAF=2 NF=2.612)
.MODEL JADJMOD NJF (BETA=4.5e-005 VTO=-1)
.MODEL DMOD D (IS=30F N=2.612)
.ENDS
*$
*
* MANUFACTURERS PART NO. = LM139   (TEXAS INSTRUMENTS)
* SUBTYPE: COMPARATOR
* THIS IS A PRE-RAD MODEL OF THE LM139 WHICH MAY BE USED
* WITH A .TEMP STATEMENT FROM -55 C TO 125 C.
* THIS MODEL MAY BE USED FOR ALL OF THE FOLLOWING DEVICES :
* LM139
* LM139J
* LM139W
* LM139A
*
*************
*
* THE FOLLOWING PARAMETERS HAVE BEEN MODELED:
* RESPONSE TIME (HL); MEAS=1US SIM=1.3US ; RESPONSE TIME (LH); MEAS=2.2US
* SIM=2US; VIO MEAS=721UV SIM=97UV; -IB MEAS=20NA SIM=15.8NA ; +IB MEAS=20NA
* SIM=17NA; IOS MEAS=132PA SIM=1.4NA; ICC+ MEAS=1.14MA SIM=1.08MA
* THIS MODEL WORKS WELL WITH ASYMMETRIC POWER SUPPLIES
*****
*
* CONNECTION:        NON-INVERTING INPUT
*                    | INVERTING INPUT
*                    | | POSITIVE POWER SUPPLY
*                    | | | NEGATIVE POWER SUPPLY
*                    | | | | OPEN COLLECTOR OUTPUT
*                    | | | | |
.SUBCKT LM139/TEMP 1 2 3 4 5
X6 3 34 LED
RE 3 35 8.4K
RS1 34 4 30.5K
Q8 7 34 35 QKI
DV1 21 1 DX
DV2 22 2 DX
Q1 9 21 7 QIN
Q2 8 22 7 QIN
Q3 9 9 4 QMO
Q4 8 9 4 QMO
Q7 11 190 19 QKI
Q6 11 8 4 QN
.MODEL QN NPN(
+         IS = 0.8F
+         BF = 250
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 7.5N
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 350N
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
RE1  3 19  8.4K
RS2 190 4 30.5K
XLED2 3 190 LED
Q5 5 11 4 QOC
.MODEL QOC NPN(
+         IS = 0.8F
+         BF = 20290
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 20N
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 1E-15
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 543.8E-9
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL QIN PNP(
+         IS = 0.8F
+         BF = 200
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 1E-15
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL QMO NPN(
+         IS = 0.8F
+         BF = 200
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 1E-15
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 807.4E-9
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL QKI PNP(
+         IS = 0.8F
+         BF = 1000
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 1E-15
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL DX D(
+         IS = 0.8F
+         RS = 0.0001
+          N = 1
+         TT = 0
+        CJO = 1E-15
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.ENDS LM139/TEMP
*
.SUBCKT LED  1      3
********** ANODE  CATHODE
D1 1 2 DX1
VL 2 3 0.8
.MODEL DX1 D(
+         IS = 0.8F
+         RS = 1
+          N = 1
+         TT = 0
+        CJO = 1E-15
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.ENDS LED
*$
* LM150 voltage regulator "macromodel" subcircuit
* created using Parts release 5.3 on 04/08/93 at 12:05
* PARTS is a MicroSim product.
*
* connections:     input
*                  |  adjustment pin
*                  |  |   output
*                  |  |   |
.SUBCKT LM150     IN ADJ OUT
*
* POSITIVE ADJUSTABLE VOLTAGE REGULATOR
*
JADJ IN ADJ ADJ JADJMOD ;ADJUSTMENT PIN CURRENT
VREF 4 ADJ 1.25
DBK IN 13 DMOD
*
* ZERO OF RIPPLE REJECTION
*
CBC 13 15 8e-010
RBC 15 5 1000
*
QPASS 13 5 OUT QPASSMOD
RB1 7 6 1
RB2 6 5 128.3
*
* CURRENT LIMITING
*
DSC 6 11 DMOD
ESC 11 OUT VALUE {11.55-0.3749*V(6,5)*V(13,5)}
*
* FOLDBACK CURRENT
*
DFB 6 12 DMOD
EFB 12 OUT VALUE {18.9-1.228*V(13,5)+0.02328*V(13,5)*V(13,5)
+ -0.374894*V(13,5)*V(6,5)}
*
EB 7 OUT 8 OUT 13.53
*
* ZERO OF OUTPUT IMPEDANCE
*
RP 9 8 100
CPZ 10 OUT 1.592e-005
*
DPU 10 OUT DMOD ;POWER-UP CLAMPLING DIODE
RZ 8 10 0.1
EP 9 OUT 4 OUT 100
RI OUT 4 100MEG
*
.MODEL QPASSMOD NPN (IS=30F BF=50 VAF=2.667 NF=2.612)
.MODEL JADJMOD NJF (BETA=5e-005 VTO=-1)
.MODEL DMOD D (IS=30F N=2.612)
.ENDS
*$
* LM196 voltage regulator "macromodel" subcircuit
* created using Parts release 5.3 on 04/08/93 at 11:33
* PARTS is a MicroSim product.
*
* connections:     input
*                  |  adjustment pin
*                  |  |   output
*                  |  |   |
.SUBCKT LM196     IN ADJ OUT
*
* POSITIVE ADJUSTABLE VOLTAGE REGULATOR
*
JADJ IN ADJ ADJ JADJMOD ;ADJUSTMENT PIN CURRENT
VREF 4 ADJ 1.25
DBK IN 13 DMOD
*
* ZERO OF RIPPLE REJECTION
*
CBC 13 15 8e-010
RBC 15 5 1000
*
QPASS 13 5 OUT QPASSMOD
RB1 7 6 1
RB2 6 5 128.3
*
* CURRENT LIMITING
*
DSC 6 11 DMOD
ESC 11 OUT VALUE {25.66-0.003981*V(6,5)*V(13,5)}
*
* FOLDBACK CURRENT
*
DFB 6 12 DMOD
EFB 12 OUT VALUE {38.46-3.533*V(13,5)+0.08855*V(13,5)*V(13,5)
+ -0.02*V(13,5)*V(6,5)}
*
EB 7 OUT 8 OUT 26.85
*
* ZERO OF OUTPUT IMPEDANCE
*
RP 9 8 100
CPZ 10 OUT 1.592e-006
*
DPU 10 OUT DMOD ;POWER-UP CLAMPLING DIODE
RZ 8 10 0.1
EP 9 OUT 4 OUT 100
RI OUT 4 100MEG
*
.MODEL QPASSMOD NPN (IS=30F BF=50 VAF=251.2 NF=1.956)
.MODEL JADJMOD NJF (BETA=5e-005 VTO=-1)
.MODEL DMOD D (IS=30F N=1.956)
.ENDS
*$
* LT1084C voltage regulator "macromodel" subcircuit
* created using Parts release 5.3 on 04/08/93 at 12:23
* PARTS is a MicroSim product.
*
* connections:     input
*                  |  adjustment pin
*                  |  |   output
*                  |  |   |
.SUBCKT LT1084C   IN ADJ OUT
*
* POSITIVE ADJUSTABLE VOLTAGE REGULATOR
*
JADJ IN ADJ ADJ JADJMOD ;ADJUSTMENT PIN CURRENT
VREF 4 ADJ 1.25
DBK IN 13 DMOD
*
* ZERO OF RIPPLE REJECTION
*
CBC 13 15 8e-010
RBC 15 5 1000
*
QPASS 13 5 OUT QPASSMOD
RB1 7 6 1
RB2 6 5 128.3
*
* CURRENT LIMITING
*
DSC 6 11 DMOD
ESC 11 OUT VALUE {17.96-0.01186*V(6,5)*V(13,5)}
*
* FOLDBACK CURRENT
*
DFB 6 12 DMOD
EFB 12 OUT VALUE {16.63+0.5959*V(13,5)-0.0801*V(13,5)*V(13,5)
+ -0.0118552*V(13,5)*V(6,5)}
*
EB 7 OUT 8 OUT 18.79
*
* ZERO OF OUTPUT IMPEDANCE
*
RP 9 8 100
CPZ 10 OUT 1.592e-005
*
DPU 10 OUT DMOD ;POWER-UP CLAMPLING DIODE
RZ 8 10 0.1
EP 9 OUT 4 OUT 100
RI OUT 4 100MEG
*
.MODEL QPASSMOD NPN (IS=30F BF=50 VAF=84.35 NF=1.373)
.MODEL JADJMOD NJF (BETA=5.5e-005 VTO=-1)
.MODEL DMOD D (IS=30F N=1.373)
.ENDS
*$
* TL783C voltage regulator "macromodel" subcircuit
* created using Parts release 5.3 on 04/08/93 at 15:09
* PARTS is a MicroSim product.
*
* connections:     input
*                  |  adjustment pin
*                  |  |   output
*                  |  |   |
.SUBCKT TL783C    IN ADJ OUT

*
* POSITIVE ADJUSTABLE VOLTAGE REGULATOR
*
JADJ IN ADJ ADJ JADJMOD ;ADJUSTMENT PIN CURRENT
VREF 4 ADJ 1.27
DBK IN 13 DMOD
*
* ZERO OF RIPPLE REJECTION
*
CBC 13 15 8e-010
RBC 15 5 1000
*
QPASS 13 5 OUT QPASSMOD
RB1 7 6 1
RB2 6 5 85.21
*
* CURRENT LIMITING
*
DSC 6 11 DMOD
ESC 11 OUT VALUE {1.96-0.01057*V(6,5)*V(13,5)}
*
* FOLDBACK CURRENT
*
DFB 6 12 DMOD
EFB 12 OUT VALUE {2.326-0.03221*V(13,5)+0.0001421*V(13,5)*V(13,5)
+ -0.02*V(13,5)*V(6,5)}
*
EB 7 OUT 8 OUT 8.069
*
* ZERO OF OUTPUT IMPEDANCE
*
RP 9 8 100
CPZ 10 OUT 1.989e-006
*
DPU 10 OUT DMOD ;POWER-UP CLAMPLING DIODE
RZ 8 10 0.1
EP 9 OUT 4 OUT 100
RI OUT 4 100MEG
*
.MODEL QPASSMOD NPN (IS=30F BF=50 VAF=94.64 NF=7.604)
.MODEL JADJMOD NJF (BETA=8.3e-005 VTO=-1)
.MODEL DMOD D (IS=30F N=7.604)
.ENDS
*$
*
*---------------------------------------------------------------------------------------

*** Voltage regulators (negative)

.SUBCKT x_LM79XX Input Output Ground PARAMS:
+       Av_feedback=1660, R1_Value=4615,
+       Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+       Rout_Value=0.01, Rreg_Value=1.2k
*
* SERIES 3-TERMINAL NEGATIVE REGULATOR
*
* Note: This regulator is based on the LM79XX series of
*       regulators (also the LM120 and LM320).  The
*       LM79XX regulators are unstable and will
*       oscillate unless a 1 uFarad solid tantalum
*       capacitor is placed on the output with an ESR
*       betweed .5 and 1.5.  This model is stable without
*       a capacitor on the output.  When performing
*       simulations a 1 uFarad capacitor should still be
*       placed on the output.  However, it it not necessary
*       to include a resistor in series with this capacitor
*       to model the ESR of the capacitor.  See the
*       comments and circuit description of the x_LM78XX
*       regulator for more information on this model.
*
* Band-gap voltage source:
*
Vbg 100 0 DC -7.4V
Sbg (100,101),(Ground,Input) Sbg1
Rbg 101 0 Rbg1 1
.MODEL Rbg1 RES (Tc1={Rbg_Tc1},Tc2={Rbg_Tc2})
Ebg (102,0),(Input,Ground) 1
Rreg 102 101 {Rreg_Value}
.MODEL Sbg1 VSWITCH (Ron=1 Roff=1MEG Von=3.7 Voff=3)
*
* Feedback stage
*
Rfb 9 8 1MEG
Cfb 8 Ground 265PF
* Eopamp 105 0 VALUE={2250*v(101,0)+Av_feedback*v(Ground,8)}
Vgainf 200 0 {Av_feedback}
Rgainf 200 0 1
Eopamp 105 0 POLY(3),(101,0),(Ground,8),(200,0) 0 2250 0 0 0 0 0 0 1
Ro 105 106 1k
D1 108 106 Dlim
D2 106 107 Dlim
.MODEL Dlim D (Vj=0.7)
Vl1 108 102 DC 1
Vl2 0 107 DC 1
*
* Quiescent current modelling
*
Gq (Ground,Input),(9,Input) 9.0E-7
R1 9 Ground {R1_Value} TC=0.001
Fl (Ground,0) Vmon 3.0E-4
*
* Output Stage
*
Q1 9 5 6 Npn1
Q2 9 6 7 Npn1 10
.MODEL Npn1 NPN (Bf=50 Is=1E-14)
* Efb 4 Ground VALUE={v(Input,Ground)+v(0,106)}
Efb 4 Ground POLY(2),(Input,Ground),(0,106) 0 1 1
Rb 4 5 1k TC=0.003
Re 6 7 2k
Rsc 7 Input 0.13 TC=1.136E-3,-7.806E-6
Rout 9 Imon {Rout_Value}
Vmon Imon Output DC 0.0
*
* Current Limit
*
Qcl1 54 52 53 Npn1
Qcl3 Input 54 5 Pnp1
.MODEL Pnp1 PNP (Bf=250 Is=1E-14)
Rcl3 5 54 1.8k
Qcl2 52 52 51 Npn1
Veset 53 Input DC 0.3v
Ibias Input 52 DC 300u
Rcl1 50 51 20k
Rcl2 51 7 115
Dz1 50 9 Dz
.MODEL Dz D (Is=0.05p Rs=3 Bv=7.11 Ibv=0.05u)
.ENDS
*$
*
*---------------------------------------------------------------LM7905C
.SUBCKT LM7905C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=1660, R1_Value=4615,
+     Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+     Rout_Value=0.01, Rreg_Value=1.2k
.ENDS
*$
*
*---------------------------------------------------------------uA7905C
.SUBCKT uA7905C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=1660, R1_Value=4615,
+     Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+     Rout_Value=0.01, Rreg_Value=1.2k
.ENDS
*$
*
*---------------------------------------------------------------LAS1805
.SUBCKT LAS1805 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=1660, R1_Value=4615,
+     Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+     Rout_Value=0.01, Rreg_Value=1.2k
.ENDS
*$
*
*---------------------------------------------------------------MC7905C
.SUBCKT MC7905C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=1660, R1_Value=4615,
+     Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+     Rout_Value=0.01, Rreg_Value=1.2k
.ENDS
*$
*
*---------------------------------------------------------------SG7905C
.SUBCKT SG7905C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=1660, R1_Value=4615,
+     Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+     Rout_Value=0.01, Rreg_Value=1.2k
.ENDS
*$
*
*---------------------------------------------------------------UC7905C
.SUBCKT UC7905C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=1660, R1_Value=4615,
+     Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+     Rout_Value=0.01, Rreg_Value=1.2k
.ENDS
*$
*
*---------------------------------------------------------------LM7912C
.SUBCKT LM7912C INPUT OUTPUT GROUND



x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=9.1k
.ENDS
*$
*
*---------------------------------------------------------------uA7912C
.SUBCKT uA7912C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=9.1k
.ENDS
*$
*
*---------------------------------------------------------------
.SUBCKT LAS1812 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=9.1k
.ENDS
*$
*
*---------------------------------------------------------------MC7912C
.SUBCKT MC7912C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=9.1k
.ENDS
*$
*
*---------------------------------------------------------------SG7912C
.SUBCKT SG7912C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=9.1k
.ENDS
*$
*
*---------------------------------------------------------------UC7912C
.SUBCKT UC7912C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=9.1k
.ENDS
*$
*
*---------------------------------------------------------------LM7915C
.SUBCKT LM7915C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=555, R1_Value=13845,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=11.3k
.ENDS
*$
*
*---------------------------------------------------------------uA7915C
.SUBCKT uA7915C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=555, R1_Value=13845,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=11.3k
.ENDS
*$
*
*---------------------------------------------------------------LAS1815
.SUBCKT LAS1815 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=555, R1_Value=13845,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=11.3k
.ENDS
*$
*
*---------------------------------------------------------------MC7915C
.SUBCKT MC7915C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=555, R1_Value=13845,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=11.3k
.ENDS
*$
*
* MANUFACTURERS PART NO.= SG7915AIG
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMP. DEPENDENT MODEL OF THE SG7915
* REGULATOR
*
*------------------------------------------------------------------------------
*
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT.  IT
* INCLUDES POWER-UP AND POWER-DOWN EFFECTS.
* IT IS NECESSARY TO SET ITL1=300 ITL2=300 WITH THE
* .OPTIONS COMMAND FOR 100% CONVERGENCE.  THESE SETTINGS DETERMINE THE
* NUMBER OF ITERATIONS ALLOWED FOR THE CALCULATION OF THE DC AND BIAS PT
* VALUES WHEN THE STARTING POINT IS CONSIDERED "BLIND" OR AN "EDUCATED
* GUESS".   OTHER SETTINGS MAY WORK, BUT HAVE NOT BEEN TESTED YET.
*
*
.SUBCKT SG7915  1 2 3 100
*               |       |   |    |
*             GND(PIN)  |   |    |
*                      OUT  |    |
*                          IN    |
*                              ZERO REFERENCE(EXTERNAL GND)
*** VOLTAGE REFERENCE SECTION ***
LZR 4 1 IND1 0.2079M
.MODEL IND1 IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 0.021188
+        TC2 = 3.9548E-4
+ )
DZR  29 4 DZR
.MODEL DZR D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 2.7117
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -2.4708E-5
+       TBV2 = 3.1346E-7
+       TRS1 = 0
+       TRS2 = 0
+ )
RZR 29 4 1MEG
RR   29 15 5.8475 TC=0.013783, 2.0804E-4
RQ   15 22 42072.4191 TC=0.007522, 1.3907E-4
D1   3 22 D1
.MODEL D1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 2
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -0.004583
+       TBV2 = 2.08333E-5
+       TRS1 = 0
+       TRS2 = 0
+ )
****
FQ 1 3 POLY(3) VQ1 VQ2 VQ3 0 1 1 -1
*** ERROR AMPLIFIER SECTION ***
EA 9 3 5 15 600
RO 6 9 200
D+ 6 20 DC
E+ 20 21 1 3 1
V+ 21 3 -1
D- 19 6 DC
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
V- 19 3 DC 1
***
RP 6 7 1
CP 7 3 1U
*** QUIESCENT CURRENT SECTION ***
EQ1 23 100 TABLE {V(1,3)} (2,100) (6.5,4.5)
VQ1 23 24 DC 0
RQ1 24 100 2251.1256 TC=0.004046, 1.1071E-5
EQ2 25 100 TABLE {V(1,3)} (6.5,0) (16,9.5)
VQ2 25 26 DC 0
RQ2 26 100 5757.81 TC=0.008862, 5.369E-5
EQ3 27 100 TABLE {V(1,3)} (16,0) (16.5,0.5)
VQ3 27 28 DC 0
RQ3 28 100 155.4 TC=0.005318, 1.2798E-5
***
GB 1 8 1 15 4M
GCOMP 3 1 1 15 4M
DB 8 18 DB
.MODEL DB D(
+         IS = 1E-14
+         RS = 0.1
+          N = 0.1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
EB 18 3 7 3 1
RB 8 10 10
*** CURRENT LIMIT AND FOLDBACK CURRENT SECTION ***
QL 1 14 14 QTEMP
.MODEL QTEMP NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
RFB 12 14 46.8663K TC=0.003476, -3.2976E-6
DZFB 13 12 DZFB
.MODEL DZFB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 7.8523
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -0.001336
+       TBV2 = 9.3921E-6
+       TRS1 = 0
+       TRS2 = 0
+ )
QCL 10 13 3 QMOD
RBCL 13 17 1K
RCL 17 3 0.2175 TC=6.659E-4, 7.318E-6
***
RBC  11 14 1762
CBC  10 11 1N
*** OUTPUT TRANSISTOR ***
QP 16 10 17 QMOD
.MODEL QMOD NPN(
+         IS = 1E-14
+         BF = 70000
+         NF = 1
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
DDO  14 30 DDO
.MODEL DDO D(
+         IS = 1E-14
+         RS = 0
+          N = 1.0876
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
RDDO 30 16 0.1
R23 1 5 2.69K
R22 5 14 12.5K
ROUT 14 2 0.0891 TC=0.003976, -2.8869E-5
DDIS 3 14 DDIS
.MODEL DDIS D(
+         IS = 1E-12
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS SG7915
*$
*
*---------------------------------------------------------------SG7915C
.SUBCKT SG7915C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=555, R1_Value=13845,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=11.3k
.ENDS
*$
*
*---------------------------------------------------------------UC7915C
.SUBCKT UC7915C Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=555, R1_Value=13845,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.01, Rreg_Value=11.3k
.ENDS
*$
*
*---------------------------------------------------------------LM120K-5
.SUBCKT LM120K-5 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=1660, R1_Value=4615,
+     Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+     Rout_Value=0.03, Rreg_Value=1.2k
.ENDS
*$
*
*---------------------------------------------------------------LM120K-12
.SUBCKT LM120K-12 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.03, Rreg_Value=9.1k
.ENDS
*$
*
*---------------------------------------------------------------LM120K-15
.SUBCKT LM120K-15 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=555, R1_Value=13845,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.03, Rreg_Value=11.3k
.ENDS
*$
*
*---------------------------------------------------------------LM320K-5
.SUBCKT LM320K-5 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=1660, R1_Value=4615,
+     Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+     Rout_Value=0.03, Rreg_Value=1.2k
.ENDS
*$
*
*---------------------------------------------------------------LM320K-12
.SUBCKT LM320K-12 Input  Output  Ground
x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.03, Rreg_Value=9.1k
.ENDS
*$
*
*---------------------------------------------------------------LM320K-15
.SUBCKT LM320K-15 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=555, R1_Value=13845,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.03, Rreg_Value=11.3k
.ENDS
*$
*
*---------------------------------------------------------------LM320T-5
.SUBCKT LM320T-5 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=1660, R1_Value=4615,
+     Rbg_Tc1=8.13E-5, Rbg_Tc2=0.0,
+     Rout_Value=0.03, Rreg_Value=1.2k
.ENDS
*$
*
*---------------------------------------------------------------LM320T-12
.SUBCKT LM320T-12 Input Output Ground
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=694, R1_Value=11076,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.03, Rreg_Value=9.1k
.ENDS
*$
*
*---------------------------------------------------------------LM320T-15
.SUBCKT LM320T-15 nput Output round
   x1 Input Output Ground x_LM79XX PARAMS:
+     Av_feedback=555, R1_Value=13845,
+     Rbg_Tc1=-9.50E-7, Rbg_Tc2=-6.53E-7,
+     Rout_Value=0.03, Rreg_Value=11.3k
.ENDS
*$
*------------------------------------------------------------------------

*** Precision voltage regulators

*---------------------------------------------------------------LM723
* connections:   current limit
*                | current sense
*                | | inverting input
*                | | | non-inverting input
*                | | | | Vref
*                | | | | | Vcc-
*                | | | | | | Vz
*                | | | | | | | Vout
*                | | | | | | | |  Vc
*                | | | | | | | |  |  Vcc+
*                | | | | | | | |  |  |  frequency compensation
*                | | | | | | | |  |  |  |
.SUBCKT LM723    2 3 4 5 6 7 9 10 11 12 13
*
* Note: This model is based on the National LM723 voltage
*       regulator.  All characterization is from data sheet
*       information.  The pin configuration corresponds to
*       the dual-in-line package.  Therefore, it includes
*       an internal 6.2 volt zener diode between Vout and Vz
*       In the model, GIee & GIcc adjust the short circuit
*       current limit and the standby current.  Rsb and the
*       temperature coefficient on RIee also affect the
*       standby current.  Bf and the transresistance term
*       on HVref adjust the low frequency output impedence
*       and the load regulation.  Rlnreg controls the line
*       regulation and ripple rejection.  Rref and its
*       temperature coefficient determine the average
*       temperature coefficient with respect to the output
*       voltage.
*
* Standby Current Correction
*
Rsb 12 7 300k
*
* Error Amplifier
*
Rlnreg 12 13 4meg
* Icc 12 13 DC 583ua
* Iee 20  7 DC 1166ua
Iee   0 24 1166ua
RIee 24 0 1 TC=4E-3
GIee (20,7),(24,0) 1.0
GIcc (12,13),(24,0) 0.5
Q5 12 5 20 Npn1
Q4 13 4 20 Npn1
*
* Voltage Reference
*
HVref 22 7 POLY(1) Vmon 7.15 0.0
Rref 22 6 15ohm TC=0.01
*
* Output Stage
*
Q1 12 13 21 Npn1
Q2 11 21 23 Npn1
Vmon 23 10 DC 0.0
Re 21 10 15k
.MODEL Npn1 NPN (Bf=55 Is=1E-14)
*
* Frequency Compensation, Current Limit, Current Sense
*
Q3 13 2 3 Npn1
R2 2  7 1.0e12
R3 3  7 1.0e12
*
* Zener Diode (6.2V) to pin 9
*
Dz 9 10 Dz
Rz 9  7 1.0e12
.MODEL Dz D (Is=0.05p Rs=4 Bv=5.79 Ibv=0.05u)
*
.ENDS
*$
*
*---------------------------------------------------------------uA723M
.SUBCKT uA723M 2 3 4 5 6 7 9 10 11 12 13
*
   x1 2 3 4 5 6 7 9 10 11 12 13 LM723
*
* the uA723M is identical to the LM723
*
.ENDS
*$
*
*---------------------------------------------------------------LM723C
.SUBCKT LM723C 2 3 4 5 6 7 9 10 11 12 13
*
   x1 2 3 4 5 6 7 9 10 11 12 13 LM723
*
* the LM723C is identical to the LM723,
* but with a more limited temperature range
*
.ENDS
*$
*
*---------------------------------------------------------------uA723C
.SUBCKT uA723C 2 3 4 5 6 7 9 10 11 12 13
*
   x1 2 3 4 5 6 7 9 10 11 12 13 LM723
*
* the uA723C is identical to the LM723,
* but with a more limited temperature range
*
.ENDS
*$
*
* MANUFACTURERS PART NO. = UA723  (FAIRCHILD)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD ROOM TEMPERATURE MODEL.
*
* * CONNECTIONS:    CURRENT SENSE
*                   | INVERTING INPUT
*                   | | NON-INVERTING INPUT
*                   | | | VREF
*                   | | | | VCC-
*                   | | | | | VOUT
*                   | | | | | | VC
*                   | | | | | | |  VCC+
*                   | | | | | | |  |  FREQUENCY COMPENSATION
*                   | | | | | | |  |  | CURRENT LIMITING
*                   | | | | | | |  |  | |
.SUBCKT UA723/27C   1 2 3 4 5 6 7  8  9 10
*
DZ1 13 8 DZ1
.MODEL DZ1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.2
+        IBV = .001
+ )
RQ 12 13 288K
R1 12 5 5.875MEG
DREF 11 12 DREF
.MODEL DREF D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 7
+        IBV = .001
+ )
RR1 11 5 700K
RR2 18 5 600
LREF 18 11 2M
RLREF 18 11 100MEG
FLOADR 5 12 VSENSE 89.35U
GQ1 8 4 12 5 0.2857M
EREF 4 5 12 5 1
RIN 2 3 100K
GQ2 8 17 4 5 0.0249M
DB 17 19 DB
.MODEL DB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
ROUT 19 14 5
EA 14 5 3 2 600
DCLOW 5 19 DCLOW
.MODEL DCLOW D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
EC 20 5 8 5 1
DCHIGH 19 20 DCHIGH
.MODEL DCHIGH D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
RB1 17 9 10
RB2 9 21 10
QL4 8 21 16 QPASS
QL5 7 16 15 QPASS
.MODEL QPASS NPN (
+         IS = 1E-16
+         BF = 50
+         NF = 1
+        VAF = 100
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
VSENSE 15 6 DC 0
RE 16 15 15K
QLIMIT 9 10 1 QLIMIT
.MODEL QLIMIT NPN  (
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.ENDS UA723/27C
*$
*
* MANUFACTURERS PART NO. = UA723  (FAIRCHILD)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT MODEL.
*
*------------------------------------------------------------------------------
*
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT. IT
* INCLUDES POWER-UP AND POWER-DOWN EFFECTS.  IT IS NECESSARY TO SET
* ITL1=300 ITL2=300 WITH THE .OPTIONS COMMAND FOR 100% CONVERGENCE. THESE
* SETTINGS DETERMINE THE NUMBER OF ITERATIONS ALLOWED FOR THE
* CALCULATION OF THE DC AND BIAS PT VALUES WHEN THE STARTING POINT IS
* CONSIDERED "BLIND" OR AN "EDUCATED GUESS". OTHER SETTINGS MAY WORK, BUT
* HAVE NOT BEEN TESTED YET.
*
*
* CONNECTIONS:        CURRENT SENSE
*                     | INVERTING INPUT
*                     | | NON-INVERTING INPUT
*                     | | | VREF
*                     | | | | VCC-
*                     | | | | | VOUT
*                     | | | | | | VC
*                     | | | | | | |  VCC+
*                     | | | | | | |  |  FREQUENCY COMPENSATION
*                     | | | | | | |  |  |  CURRENT LIMITING
*                     | | | | | | |  |  | |   GND(REFERENCE)
.SUBCKT UA723/TEMP    1 2 3 4 5 6 7  8  9 10  99
*
*** REFERENCE SECTION ***
DZ1 13 8 DZ1
.MODEL DZ1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1
+        IBV = .001
+ )
RQ 40 13 237.273K TC=2.7132E-3, 6.8655E-6
DZR 11 40 DZR
.MODEL DZR D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 6.9504
+        IBV = .001
+ )
RZR 11 40 1MEG
RR1 11 500 100.1936 TC=6.4819E-3, -5.0748E-6
LR 500 5 LR 1.139M
.MODEL LR IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 8.1788E-3
+        TC2 = 2.1531E-5
+ )
RR2 500 5 15K
CR 11 1000 3P
RCR 1000 5 10
*** CURRENT SOURCE ***
GQ1 8 4 POLY(2) (4,5) (10000,99) 0 0.2832M 0 0 -2.2853E-7 0 0 0 -1.8472E-10
GQ2 8 17 4 5 0.08M
ER 4 5 40 5 1
RIN 2 3000 100K
HLDR 3 3000 POLY(2) VLDR VT 0 35.2M 0 0 -4.6889E-5 0 0 0 9.03892E-6
*** FREQUENCY COMP ERROR AMPLIFIER ***
DB 17 19 DB
.MODEL DB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
RO 19 14 500
EA 14 5 3000 2 600
D- 22 19 DC
V- 22 5 DC 1
E+ 23 5 8 5 1
D+ 19 20 DC
V+ 20 23 DC -1.6
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
*** TEMPERATURE CHANGE CIRCUITRY ***
RT1 10000 10001 100.00001 TC=0.01
RT2 10001 99 -100.00001
IT 99 10000 DC 1
GT 99 30000 10000 99 1
VT 30000 30001 DC 0
RT3 30001 99 1
*** SERIES PASS AMPLIFIER ***
RB1 17 9 10
RB2 9 21 10
QP1 8 21 16 QPASS1
QP2 7 16 15 QPASS2
.MODEL QPASS1 NPN (
+         IS = 1E-20
+         BF = 50
+         NF = 1.0188
+        VAF = 50
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
.MODEL QPASS2 NPN (
+         IS = 1E-20
+         BF = 50
+         NF = 1.0188
+        VAF = 50
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
CBC1 8 800 1P
RCBC1 21 800 10
CBC2 7 160 1P
RCBC2 160 16 10
*** CURRENT LIMITING BLOCK ***
VLDR 15 6 DC 0
QL 9 125 1 QLIMIT
.MODEL QLIMIT NPN(
+         IS = 1E-20
+         BF = 100
+         NF = 1.3464
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
ESC 10 125 POLY(1) (10000,99) 0 -0.002738 -6.274E-5
DDIS1 6 8 DDIS
.MODEL DDIS D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS UA723/TEMP
*$
*
*---------------------------------------------------------------MC1723C
.SUBCKT MC1723C 2 3 4 5 6 7 9 10 11 12 13
*
   x1 2 3 4 5 6 7 9 10 11 12 13 LM723
*
* the MC1723C is identical to the LM723,
* but with a more limited temperature range
*
.ENDS
*$
*
*---------------------------------------------------------------CA723
.SUBCKT CA723 2 3 4 5 6 7 9 10 11 12 13
*
   x1 2 3 4 5 6 7 9 10 11 12 13 LM723
*
* the CA723 is identical to the LM723,
* but with a more limited temperature range
*
.ENDS
*$
*
* MANUFACTURERS PART NO. = CA3085BT/3  (RCA)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT MODEL OF THE CA3085.
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT. IT
* INCLUDES POWER-UP AND POWER-DOWN EFFECTS.
* IT IS NECESSARY TO SET ITL1=300 ITL2=300 WITH THE .OPTIONS COMMAND FOR
*.100% CONVERGENCE. THESE SETTINGS DETERMINE THE NUMBER OF ITERATIONS
* ALLOWED FOR THE CALCULATION OF THE DC AND BIAS PT VALUES WHEN THE STARTING
* POINT IS CONSIDERED "BLIND" OR AN "EDUCATED GUESS". OTHER SETTINGS MAY
* WORK, BUT HAVE NOT BEEN TESTED YET.
*
*
*
.SUBCKT CA3085  1    2  3  4 5 6 7 8 100
*             VOUT   |  |  | | | | |  |
*                    CB |  | | | | |  |
*                      VIN | | | | |  |
*                         V- | | | |  |
*                         VREF | | |  |
*                            IN- | |  |
*                             COMP |  |
*                              CLIMIT |
*                   GND(REFERENCE)
*
*** REFERENCE SECTION ***
D1 3 9 DMOD
DZB 10 9 DZB
.MODEL DZB D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.9
+        IBV = .001
+ )
RQ 10 11 34.034K TC=1.7516E-3,2.7249E-6
DZR 13 11 DZR
.MODEL DZR D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.637
+        IBV = .001
+ )
LR 14 4 IND1 0.2028M
.MODEL IND1 IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 2.2862E-3
+        TC2 = 1.0471E-5
+ )
RR1 13 14 29.3092 TC=8.4331E-4,-7.3654E-5
D2 11 12 DMOD
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
RR2 11 4 43.316K
RR3 12 4 15.853K
ER 5 4 11 4 1
VLDR 22 1 DC 0
HLDR 15 6 POLY(2) VLDR VT 0 -0.0436 0 0 0.002734 0 0 0 -2.293E-5
*** CURRENT SOURCE ***
GB1 3 5 POLY(2),(12,4),(10000,100) 0 .8999M 0 0 3.6889E-6 0 0 0 -3.1779E-8
GB2 3 7 12 4 2M
*** FREQUENCY COMP ERROR AMPLIFIER ***
RIN 5 15 1MEG
DL 7 17 DL
.MODEL DL D(
+         IS = 1E-14
+         RS = 0
+          N = 0.1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
ED 18 4 5 15 10000
E+ 16 4 9 4 1
D+ 17 160 DMOD
V+ 160 16 DC -1
DC- 40 17 DMOD
V- 40 4 DC 1
*** TEMPERATURE CHANGE CIRCUITRY ***
RT1 10000 10001 100.00001 TC=0.01
RT2 10001 100 -100
IT 100 10000 DC 1
GT 100 30000 10000 0 1
VT 30000 30001 DC 0
RT3 30001 100 1
RO 17 18 5
*** SERIES PASS AMPLIFIER ***
RB 7 20 10
QP2 3 20 21 QMOD1
QP1 2 21 22 QMOD1
.MODEL QMOD1 NPN (
+         IS = 1E-16
+         BF = 50
+         NF = 1.25
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
*** CURRENT LIMITING BLOCK ***
R5 3 2 500
RB15 200 1 1.5K
QL 7 19 8 QLIMIT
.MODEL QLIMIT NPN(
+         IS = 1E-14
+         BF = 100
+         NF = 1.0666
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
EL 19 200 POLY(1),(10000,100) 0 -6.7125E-4 5.0625E-6
DDIS 1 3 DDIS
.MODEL DDIS D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS CA3085
*$
*
* MANUFACTURERS PART NO. = CA3085BT/3  (RCA)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD ROOM TEMPERATURE MODEL.
*
******
*---------------------------------------------------------------------------
* PLEASE NOTE THE FOLLOWING:
*
* 1) THIS MODEL IS TO BE USED FOR ROOM TEMPERATURE SIMULATIONS.  THE
*    SPICE TEMPERATURE CORRECTIONS WILL NOT WORK.
* 2) FOR FURTHER DETAILS AND THE MODEL DERIVATION, SEE
*    "CA3085, LM7805, LM7812, LM7905, LM137 MACROMODEL DEVELOPMENT"
*    BY G. M. WIERZBA.
*
.SUBCKT CA3085/25C 1 2 3 4 5 6 7 8
*            VOUT | | | | | | |
*                CB | | | | | |
*                 VIN | | | | |
*                    V- | | | |
*                    VREF | | |
*                       IN- | |
*                        COMP |
*                        CLIMIT
*
*
DTEST 3 300 DMOD
DZB 202 300 DZ3
.MODEL DZ3 D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 0.4
+        IBV = .001
+ )
R1 202 200 33.844K
DZR 203 200 DZ1
.MODEL DZ1 D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.605
+        IBV = .001
+ )
RR 203 4 18.2
D2 200 201 DMOD
.MODEL DMOD D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
R2 200 4 26.592K
R3 201 4 20.39035K
GBIAS1 3 5 201 4 2.9M
ER 5 4 200 4 1
RIN 5 6 0.1MEG
GBIAS2 3 7 201 4 150U
DLIMIT1 7 10 DMOD1
.MODEL DMOD1 D(
+         IS = 1E-14
+         RS = 0
+          N = 0.1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
CDLIMIT 7 10 1U
EDIFF 100 4 5 6 0.1MEG
ROUT 10 100 5
ECLAMP1 22 4 202 4 1
DCLAMP1 10 22 DMOD
DCLAMP2 4 10 DMOD1
RB 7 12 3K
CBC 12 20 0.25U
RBC 20 19 1.5K
QPASS 19 12 1000 QMOD1
RZO 1000 1 3.8
.MODEL QMOD1 NPN (
+         IS = 1E-14
+         BF = 1000
+         NF = 1
+        VAF = 50
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
DD02 2 18 DMOD2
DD01 18 19 DMOD2
.MODEL DMOD2 D(
+         IS = 1E-14
+         RS = 0
+          N = 1.3734
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
R5 3 2 500
RB15 13 1 1.5K
QLIMIT 24 13 8 QMOD2
DB 7 24 DB
.MODEL DB D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.MODEL QMOD2 NPN (
+         IS = 1E-14
+         BF = 100
+         NF = 1.1890
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.ENDS CA3085/25C
*$
*
* MANUFACTURERS PART NO. = LM137HVH  (NATIONAL SEMICONDUCTOR)
* SUBTYPE: REGULATOR
*
* THIS FILE CONTAINS A PRE-RAD MODEL AT 27 C OF THE  LM137HVH THAT WAS
* DEVELOPED UNDER THE GUIDANCE OF GREGORY M. WIERZBA AT
* MICHIGAN STATE UNIVERSITY.
*
* PLEASE NOTE THE FOLLOWING:
*
*   1) THIS MODEL IS TO BE USED FOR ROOM TEMPERATURE SIMULATIONS. THE BUILT-
*       IN  SPICE TEMPERATURE CORRECTIONS WILL NOT WORK.
*   2) RIPPLE REJECTION, OUTPUT IMPEDANCE, LINE TRANSIENT, AND LOAD
*       TRANSIENT RESPONSE ARE MODELED BASED ON LABORATORY
*       MEASUREMENTS.  THE CORRELATION IS QUITE GOOD. THE SIMULATION VALUES
*       ARE WITHIN THE PRODUCT SPEC LIMITS.
*   3) CURRENT LIMITING AND ADJUSTMENT CURRENT BASED ON DATA SHEET
*       INFORMATION ARE MODELED ACCURATELY.
*   4) DROPOUT AND POWER UP CHARACTERISTICS HAVE NOT BEEN DEVELOPED YET
*       IN THIS  MODEL.
*   5) FOR FURTHER DETAILS AND THE MODEL DERIVATION, OBTAIN A COPY OF
*      "CA3085,  LM7805, LM7812, LM7905, LM137 MACROMODEL DEVELOPMENT" BY G. M.
*        WIERZBA  DATED 3/25/91.
*
*
*
.SUBCKT LM137HVH  1  2  3
*                IN  |  |
*                   OUT |
*                      ADJ
*
VREF   12  4  DC 1.25
EREG   3  12  1  2  0.0001981
IBIAS  4  1  DC 65U
RIN    4  20 100MEG
E1     5  1  20  4  600
R1     5  6  1561
RPZ    6  11  0.01
C1     11 1  1U
E2     7  1  6  1  1
RB1    7  17  25
RB2    17  8  50
DLIMIT 17  18  DMOD
ELIMIT 18  1  POLY (1)  (2,1) .24  -0.0024
DFLDBCK 17  19   DMOD
EFLDBCK  19  1  POLY(1)  (2,1)  1.0611 -0.0912  0.0026  -2.5E-5
CBC     8  9  1U
RBC     9  20  1561
QPASS   20  8  1  QMOD
RBOND   20  2  0.0063
.MODEL QMOD NPN(
+         IS = 1E-16
+         BF = 500
+         NF = 1
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL DMOD D(
+         IS = 1E-15.9
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.ENDS LM137HVH
*$
*
* MANUFACTURERS PART # = F78M12HM
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A TEMPERATURE DEPENDENT MODEL OF THE F78M12
* REGULATOR.
*
*
*------------------------------------------------------------------------------
*
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP STATEMENT.  IT
* INCLUDES POWER-UP AND POWER-DOWN EFFECTS.
* IT IS NECESSARY TO SET ITL1=300 ITL2=300 WITH THE .OPTIONS COMMAND FOR
* 100%  CONVERGENCE.  THESE SETTINGS DETERMINE THE NUMBER OF ITERATIONS
* ALLOWED FOR  THE CALCULATION OF THE DC AND BIAS PT VALUES WHEN THE
* STARTING POINT IS  CONSIDERED "BLIND" OR AN "EDUCATED GUESS".
* OTHER SETTINGS MAY WORK, BUT HAVE NOT BEEN TESTED YET.
*
.SUBCKT F78M12  1  2   3
*               |  |   |
*              IN  |   |
*                 OUT  |
*                     GND
*
*** VOLTAGE REFERENCE AND BIAS CURRENT SECTION ***
DZ1  4 1 DZ1
.MODEL DZ1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 0.75
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -0.003611
+       TBV2 = 6.9444E-5
+       TRS1 = 0
+       TRS2 = 0
+ )
RQ   4 17 86343.84 TC=5.3597E-4, 5.0408E-5
RR   17 18 5.2447 TC=0.005772, 6.2073E-5
DZR   16 18 DR
.MODEL DR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.2588
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 3.82E-5
+       TBV2 = -8.5068E-7
+       TRS1 = 0
+       TRS2 = 0
+ )
RZ 16 18 1MEG
L1 16 3 IND1 0.3573M
.MODEL IND1 IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 0.001123
+        TC2 = 6.8566E-5
+ )
*** ERROR AMPLIFIER SECTION ***
EA 22 3 17 15 300
ROUT 22 6 10
D- 3 6 DCLAMP
D+ 6 19 DCLAMP
.MODEL DCLAMP D  (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
V+ 19 23 DC -1
E+ 23 3 1 3 1
RP 6 7 500
CP 7 3 CAP1 0.1U
.MODEL CAP1 CAP(
+          C = 1
+        VC1 = 0
+        VC2 = 0
+        TC1 = -0.002
+        TC2 = 1E-4
+ )
*** QUIESCENT CURRENT ***
GB 1 9 17 3 0.4944M
RQUIES 12 3 10572.61 TC=0.013985, 1.28953E-4
*** SHORT CIRCUIT AND FOLDBACK CURRENT ***
DBL 9 8 DBL
.MODEL DBL D(
+         IS = 1E-4
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 0
+        XTI = 0
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
EB 8 3 7 3 2
RC 1 14 0.2
DC 14 13 DC
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1.6339
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
RB 9 11 100
QP 13 11 5 QP
.MODEL QP NPN(
+         IS = 1E-12
+         BF = 70K
+         NF = 1
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
DCL 9 10 DCL
.MODEL DCL D(
+         IS = 1E-4
+         RS = 0
+          N = 2
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
QCL 10 20 12 QCL
.MODEL QCL NPN(
+         IS = 1E-16
+         BF = 100
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
RSC 5 12 0.6936 TC=0.00131, 1.2433E-5
RBCL 20 5 200
RFB 1 21 6.17043K TC=0.001143, -1.081421E-5
DZFB 20 21 DZFB
.MODEL DZFB D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 14.79
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.01
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -1.78236E-4
+       TBV2 = 4.2164E-6
+       TRS1 = 0
+       TRS2 = 0
+ )
R24 15 3 600
R23 12 15 5160
*** OUTPUT RESISTANCE ***
RO 12 2 0.02 TC=-8.3333E-4, -4.1667E-5
DDIS 2 1 DMOD
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 0.7
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS F78M12
*$
*
*---------------------------------------------------------------RC723
.SUBCKT RC723 2 3 4 5 6 7 9 10 11 12 13
*
   x1 2 3 4 5 6 7 9 10 11 12 13 LM723
*
* the RC723 is identical to the LM723,
* but with a more limited temperature range
*
.ENDS
*$
*
* MANUFACTURERS PART NO.= SG137A   (SILICON GENERAL)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD TEMPERATURE DEPENDENT MACROMODEL OF THE
* SG137A.
*
* PLEASE NOTE THE FOLLOWING:
*
* THIS MODEL CAN BE USED FROM -55 C TO 125 C WITH THE .TEMP
* STATEMENT.  IT INCLUDES POWER-UP AND POWER-DOWN EFFECTS.    IT IS
* NECESSARY TO SET ITL1=300  ITL2=300 WITH THE .OPTIONS COMMAND FOR 100%
* CONVERGENCE.  THESE  SETTINGS DETERMINE THE NUMBER OF ITERATIONS
* ALLOW FOR THE  CALCULATION OF THE DC AND BIAS PT VALUES WHEN THE
* STARTING POINT  IS CONSIDERED "BLIND" OR AN "EDUCATED GUESS".
* OTHER SETTINGS MAY WORK, BUT HAVE NOT BEEN TESTED YET.
*
* RIPPLE REJECTION, OUTPUT IMPEDANCE, QUIESCENT CURRENT, LINE
* TRANSIENT, DROPOUT, AND LOAD TRANSIENT RESPONSE ARE MODELED BASED
* ON LABORATORY MEASUREMENTS.  THE CORRELATION IS QUITE GOOD.
* CURRENT LIMITING AND ADJUSTMENT CURRENT BASED ON DATA SHEET
* INFORMATION ARE MODELED ACCURATELY.
*
*
*------------------------------------------------------------------
*
*
*
.SUBCKT SG137   1  2   3   100
*               |  |   |    |
*              ADJ |   |    |
*                 OUT  |    |
*                     IN    |
*                          GND(REFERNCE)
*** VOLTAGE REFERENCE SECTION ***
LR 1 4 IND1 0.2709
.MODEL IND1 IND(
+          L = 1
+        IL1 = 0
+        IL2 = 0
+        TC1 = 7.8864E-4
+        TC2 = -2.8391E-5
+ )
RR 4 5 98.2994 TC=-0.0063, 6.2251E-5
CR 1 6 3P
RCR 6 7 150K
DZR 7 5 DZR
.MODEL DZR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0.1P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.25
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.0001
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 2.2444E-6
+       TBV2 = 6.5556E-8
+       TRS1 = 0
+       TRS2 = 0
+ )
RZR 7 5 1MEG
DZ1 8 7 DZ1
.MODEL DZ1 D(
+         IS = 1E-14
+         RS = 1
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 0.0001
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = -0.002847
+       TBV2 = 3.4722E-6
+       TRS1 = 0
+       TRS2 = 0
+ )
RQ 8 3 1.7546MEG TC=4.5212E-4,5.6515E-6
*** QUIESCENT CURRENT SECTION ***
FQ  1 3 VQ1 0.0625M
EQ1 24 100 1 7 1
VQ1 24 25 DC 0
RQ1 25 100 1 TC=-3.9528E-4,-1.1597E-5
*** ERROR AMPLIFIER ***
RIN 7 23 100K
E1  11 3 23 7 600
ROE1 9 11 10
D+ 9 13 DC
V+ 14 3 -1
E+ 13 14 1 3 1
.MODEL DC D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 10P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
D- 12 9 DC
V- 12 3 DC 1
RP 9 10 151
CP 10 3 0.01U
E2 15 3 10 3 1
***
RB1 15 16 50
RB2 16 19 500 TC=-1.9327E-4,3.3434E-6
*** SHORT CIRCUIT AND FOLDBACK CURRENT SECTION ***
DSC 16 17 DMOD
ESC 17 3 POLY(1),(2,3) 2.447 -0.01
DFB 16 18 DMOD
EFB 18 3 POLY(1),(2,3) 12.5955 -1.2275 0.0457 -5.9169E-4
***
QP 20 19 3 QMOD
.MODEL QMOD NPN(
+         IS = 1E-14
+         BF = 500
+         NF = 1
+        VAF = 9.9999E+13
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         NK = .5
+        ISS = 0
+         NS = 1
+        QCO = 0
+        RCO = 0
+         VO = 10
+      GAMMA = 1E-11
+       TRE1 = 0
+       TRE2 = 0
+       TRB1 = 0
+       TRB2 = 0
+       TRM1 = 0
+       TRM2 = 0
+       TRC1 = 0
+       TRC2 = 0
+ )
*** DROPOUT VOLTAGE SECTION ***
RDO 23 22 0.1
DDO1 22 21 DDO
DDO2 21 20 DDO
.MODEL DDO D(
+         IS = 1E-14
+         RS = 0
+          N = 0.9687
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
***
RO 23 2 0.0017 TC=-0.07894, 0.001136
DDIS 3 23 DDIS
.MODEL DDIS D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1PF
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = 1E-10
+        ISR = 0
+         NR = 2
+        IKF = 9.9999E+13
+        NBV = 1
+       IBVL = 0
+       NBVL = 1
+       TIKF = 0
+       TBV1 = 0
+       TBV2 = 0
+       TRS1 = 0
+       TRS2 = 0
+ )
.ENDS SG137
*$
*
* MANUFACTURERS PART NO.= SG137A   (SILICON GENERAL)
* SUBTYPE: REGULATOR
* THIS FILE CONTAINS A PRE-RAD 27 C TEMP. MACROMODEL
*
*-------------------------------------------------------------------
*  PLEASE NOTE THE FOLLOWING:
* 1)  THIS MODEL IS TO BE USED FOR ROOM TEMPERATURE SIMULATIONS.
*     THE BUILT-IN SPICE TEMPERATURE CORRECTIONS WILL NOT WORK.
* 2)  RIPPLE REJECTION, OUTPUT IMPEDANCE, QUIESCENT CURRENT,
*     LINE TRANSIENT, AND LOAD TRANSIENT RESPONSE ARE MODELED
*     BASED ON LABORATORY MEASUREMENTS.  THE CORRELATION IS
*     QUITE GOOD.
* 3)  CURRENT LIMITING AND ADJUSTMENT CURRENT BASED ON DATA
*     SHEET INFORMATION ARE MODELED ACCURATELY.
* 4)  DROPOUT AND POWER UP CHARACTERISTICS HAVE NOT BEEN
*     DEVELOPED YET IN THIS MODEL.
* 5)  FOR FURTHER DETAILS AND THE MODEL DERIVATION, OBTAIN
*     A COPY OF "CA3085, LM7805, LM7812, LM7905, LM137 MACROMODEL
*     DEVELOPMENT" BY G. M. WIERZBA DATED 03/25/91.
*
*
*
.SUBCKT SG137/27C   1   2   3
*                   |   |   |
*                  IN   |   |
*                      OUT  |
*                          ADJ
RR     3 12 2250
DZR    13 12 DZR
.MODEL DZR D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 1.25
+        IBV = .001
+ )
RDZR   3 13 100MEG
D1     14 13 D1
.MODEL D1 D (
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 0.8
+        IBV = .001
+ )
RD1    14 1 14 MEG
GQ     4 1 3 13 0.052M
EREF   4 3 13 3 1
RIN    4 20 100MEG
E1     50 1 20 5 600
RCLAMP 5 50 10
EC     51 1 3 1 0.1
DCLAMP 51 5 DCLAMP
.MODEL DCLAMP D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
R1     5 6 156
RPZ    6 11 1000
C1     11 1 0.5U
E2     7 1 6 1 1
RB1    7 17 25
RB2    17 8 50
DLIMIT 17 18 DMOD
ELIMIT 18 1 POLY(1),(2,1) 0.24 -0.0024
DFLDBCK 17 19 DMOD
EFLDBCK 19 1 POLY(1),(2,1) 1.0611 -0.0912 0.0026 -2.5E-5
CBC    8 9 0.01U
RBC    9 23 10
QPASS  23 8 1 QMOD
RC     20 21 0.5
DC     21 22 DC
DO     22 23 DC
.MODEL DC D (
+         IS = 1E-14
+         RS = 0
+          N = 1.250
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
RO     20 2 0.00001
.MODEL QMOD NPN (
+         IS = 1E-16
+         BF = 500
+         NF = 1
+        VAF = 150
+        IKF = 9.9999E+13
+        ISE = 0
+         NE = 1.5
+         BR = 1
+         NR = 1
+        VAR = 9.9999E+13
+        IKR = 9.9999E+13
+        ISC = 0
+         NC = 2
+         RB = 0
+        IRB = 9.9999E+13
+        RBM = 0
+         RE = 0
+         RC = 0
+        CJE = 0
+        VJE = .75
+        MJE = .33
+         TF = 0
+        XTF = 0
+        VTF = 9.9999E+13
+        ITF = 0
+        PTF = 0
+        CJC = 0
+        VJC = .75
+        MJC = .33
+       XCJC = 1
+         TR = 0
+        CJS = 0
+        VJS = .75
+        MJS = 0
+        XTB = 0
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+ )
.MODEL DMOD D(
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 0
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 9.9999E+13
+        IBV = .001
+ )
.ENDS SG137/27C
*$
*
*---------------------------------------------------------------SG723C
.SUBCKT SG723C 2 3 4 5 6 7 9 10 11 12 13
*
   x1 2 3 4 5 6 7 9 10 11 12 13 LM723
*
* the SG723C is identical to the LM723,
* but with a more limited temperature range
*
.ENDS
*$
***** NE5532 Source: Texas Instruments NE5534
* C2 added to simulate compensated frequency response (Uwe Beis)

* NE5532 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING NE5534 model from Texas InstrumentsAT 12:41
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT NE5532   1 2 3 4 5
*
C1   11 12 7.703E-12
C2    6  7 23.500E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 2.893E6 -3E6 3E6 3E6 -3E6
GA    6  0 11 12 1.382E-3
GCM   0  6 10 99 13.82E-9
IEE  10  4 DC 133.0E-6
HLIM 90  0 VLIM 1K
Q1   11  2 13 QX
Q2   12  1 14 QX
R2    6  9 100.0E3
RC1   3 11 723.3
RC2   3 12 723.3
RE1  13 10 329
RE2  14 10 329
REE  10 99 1.504E6
RO1   8  5 50
RO2   7 99 25
RP    3  4 7.757E3
VB    9  0 DC 0
VC    3 53 DC 2.700
VE   54  4 DC 2.700
VLIM  7  8 DC 0
VLP  91  0 DC 38
VLN   0 92 DC 38
.MODEL DX D(IS=800.0E-18)
.MODEL QX NPN(IS=800.0E-18 BF=132)
.ENDS

*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Inc.
* Models developed and under copyright by:
* National Semiconductor, Inc.

*/////////////////////////////////////////////////////////////////////
* Legal Notice: This material is intended for free software support.
* The file may be copied, and distributed; however, reselling the
*  material is illegal

*////////////////////////////////////////////////////////////////////
* For ordering or technical information on these models, contact:
* National Semiconductor's Customer Response Center
*                 7:00 A.M.--7:00 P.M.  U.S. Central Time
*                                (800) 272-9959
* For Applications support, contact the Internet address:
*  Appshelp@galaxy.nsc.com

*//////////////////////////////////////////////////////////
*LM6132A OP-AMP MACRO-MODEL
*//////////////////////////////////////////////////////////
*
* Connections:      Non-inverting input
*                   |   Inverting input
*                   |   |   Positive power supply
*                   |   |   |   Negative power supply
*                   |   |   |   |   Output
*                   |   |   |   |   |
*                   |   |   |   |   |
.SUBCKT LM6132A/NS  1   2  99  50  28
* CAUTION:  SET .OPTIONS GMIN=1E-16 TO CORRECTLY MODEL INPUT BIAS CURRENT.
* Features:
* Operates from single supply
* Rail-to-rail output swing
* Offset voltage (max) = 6mV
* Input current = 170nA
* Slew rate = 27V/uS
* Gain-bandwidth product = 17MHZ
* Low supply current = 600uA
*
* NOTE: - This model is for a single device only and the simulated
*         supply current is for one op amp only.
*       - Noise is not modeled.
*       - Asymmetrical gain is not modeled.
*       - In the next revision, the following will be modelled
*       - Voltage dependent (Vin or Vcc) slew rate
*       - Gain/phase variation vs output Z
*
CI1 1  50 2P
CI2 2  50 2P
*
* 53Hz pole capacitor
C3 98 9 0.15N
*
C4  6  5  .493P
C5  98 15 2F
C7 98 11 20F
*
DP1 1  99 DA
DP2 50 1  DX
DP3 2  99 DB
DP4 50 2  DX
D1  9  8  DX
D2  10 9  DX
D3  15 20 DX
D4  21 15 DX
D5  26 24 DX
D6  25 27 DX
D7  22 99 DX
D8  50 22 DX
D9  0  14 DX
D10 12 0  DX
D11 11 33 DX
D12 34 11 DX
D14 31 32 DX
EH  97 98 99    49 1.0
EN  0  96 0     50 1.0
* Input offset voltage -|
EOS 7  1  POLY(1) 16 49 2M 1
EP  97 0  99    0  1.0
E1  97 19 99    15 1.0
E2  18 7  32    99 1E-3
* Sourcing load +Vs current
F1  99 0  VA2   1
* Sinking load -Vs current
F2  0  50 VA3   1
F3  13 0  VA1   1
G1  98 9  5     6  0.1
G2  98 11 9     49 1U
G3  98 15 11    49 1U
* DC CMRR
G4  98 16 POLY(2) 1 49 2 49 0 3.5E-9 3.5E-9
I1 99 4 18U
I2 99 50 319U
* Load dependent pole
L1 22 28 300N
*
* CMR lead
L2  16 17 7.95M
M1  5  2  4  99 MX
M2  6  18 4  99 MX
R3  5  50 1.20K
R4  6  50 1.20K
R5  98 9  1E7
R8  99 49 133.3K
R9  49 50 133.3K
R12 98 11 1E6
R13 98 17 1K
*
* -Rout
R16 23 24 62
* +Rout
R17 23 25 138
*
* +Isc slope control
R18 20 29 12K
* -Isc slope control
R19 21 30 12K
*
R21 98 15 1E6
R22 22 28 900
R23 32 97 100K
VA1 19 23 0V
VA2 14 13 0V
VA3 13 12 0V
V2  97 8  0.61V
V3  10 96 0.61V
V4  29 22 .21V
V5  22 30 .21V
V6  26 22 0.61V
V7  22 27 0.61V
V8 31 50 4V
V9 34 96 .34
V10 97 33 .34
*
.MODEL  DA D    (IS=110E-9)
.MODEL  DB D    (IS=113.4E-9)
.MODEL  DX D    (IS=1.0E-14)
.MODEL  MX PMOS (VTO=-.6 KP=4.2E-4 GAMMA=1.1)
.ENDS
*$
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Inc.
* Models developed and under copyright by:
* National Semiconductor, Inc.

*/////////////////////////////////////////////////////////////////////
* Legal Notice: This material is intended for free software support.
* The file may be copied, and distributed; however, reselling the
*  material is illegal

*////////////////////////////////////////////////////////////////////
* For ordering or technical information on these models, contact:
* National Semiconductor's Customer Response Center
*                 7:00 A.M.--7:00 P.M.  U.S. Central Time
*                                (800) 272-9959
* For Applications support, contact the Internet address:
*  Appshelp@galaxy.nsc.com

*//////////////////////////////////////////////////////////
*LM6132B OP-AMP MACRO-MODEL
*//////////////////////////////////////////////////////////
*
* Connections:      Non-inverting input
*                   |   Inverting input
*                   |   |   Positive power supply
*                   |   |   |   Negative power supply
*                   |   |   |   |   Output
*                   |   |   |   |   |
*                   |   |   |   |   |
.SUBCKT LM6132B/NS  1   2  99  50  28
* CAUTION:  SET .OPTIONS GMIN=1E-16 TO CORRECTLY MODEL INPUT BIAS CURRENT.
* Features:
* Operates from single supply
* Rail-to-rail output swing
* Offset voltage (max) = 6mV
* Input current = 170nA
* Slew rate = 27V/uS
* Gain-bandwidth product = 10MHZ
* Low supply current = 360uA
*
* NOTE: - This model is for a single device only and the simulated
*         supply current is for one op amp only.
*       - Noise is not modeled.
*       - Asymmetrical gain is not modeled.
*       - In the next revision, the following will be modelled
*       - Voltage dependent (Vin or Vcc) slew rate
*       - Gain/phase variation vs output Z
*
CI1 1  50 2P
CI2 2  50 2P
*
* 53Hz pole capacitor
C3 98 9 0.15N
*
C4  6  5  .493P
C5  98 15 2F
C7 98 11 20F
*
DP1 1  99 DA
DP2 50 1  DX
DP3 2  99 DB
DP4 50 2  DX
D1  9  8  DX
D2  10 9  DX
D3  15 20 DX
D4  21 15 DX
D5  26 24 DX
D6  25 27 DX
D7  22 99 DX
D8  50 22 DX
D9  0  14 DX
D10 12 0  DX
D11 11 33 DX
D12 34 11 DX
D14 31 32 DX
EH  97 98 99    49 1.0
EN  0  96 0     50 1.0
* Input offset voltage -|
EOS 7  1  POLY(1) 16 49 6M 1
EP  97 0  99    0  1.0
E1  97 19 99    15 1.0
E2  18 7  32    99 1E-3
* Sourcing load +Vs current
F1  99 0  VA2   1
* Sinking load -Vs current
F2  0  50 VA3   1
F3  13 0  VA1   1
G1  98 9  5     6  0.1
G2  98 11 9     49 1U
G3  98 15 11    49 1U
* DC CMRR
G4  98 16 POLY(2) 1 49 2 49 0 3.5E-9 3.5E-9
I1 99 4 18U
I2 99 50 319U
* Load dependent pole
L1 22 28 300N
*
* CMR lead
L2  16 17 7.95M
M1  5  2  4  99 MX
M2  6  18 4  99 MX
R3  5  50 1.20K
R4  6  50 1.20K
R5  98 9  1E7
R8  99 49 133.3K
R9  49 50 133.3K
R12 98 11 1E6
R13 98 17 1K
*
* -Rout
R16 23 24 62
* +Rout
R17 23 25 138
*
* +Isc slope control
R18 20 29 12K
* -Isc slope control
R19 21 30 12K
*
R21 98 15 1E6
R22 22 28 900
R23 32 97 100K
VA1 19 23 0V
VA2 14 13 0V
VA3 13 12 0V
V2  97 8  0.61V
V3  10 96 0.61V
V4  29 22 .21V
V5  22 30 .21V
V6  26 22 0.61V
V7  22 27 0.61V
V8 31 50 4V
V9 34 96 .34
V10 97 33 .34
*
.MODEL  DA D    (IS=110E-9)
.MODEL  DB D    (IS=113.4E-9)
.MODEL  DX D    (IS=1.0E-14)
.MODEL  MX PMOS (VTO=-.6 KP=4.2E-4 GAMMA=1.1)
.ENDS
*$

