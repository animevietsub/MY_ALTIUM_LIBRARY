*
*******************************************
*
*BZT52-C10
*
*Nexperia
*
*Voltage regulator diodes
*
*
*VZmax = 10,6V @ Iz = 5mA
*
*
*VFmax = 0,9V @ IF = 10mA
*IRmax = 200nA @ VR = 7V
*
*
*
*
*
*
*
*
*
*Package pinning does not match Spice model pinning.
*Package: SOD123
*
*Package Pin 1: cathode
*Package Pin 2: anode
*
*
*
*Extraction date (week/year): 04/2022
*Simulator: SPICE3
*
*******************************************
*#
.SUBCKT BZT52 1 2 PARAMS: Vbreak=10
R1 1 2 1E+12
D1 1 2
+ DIODE1
D2 1 2
+ DIODE2
*
*The resistor R1 and the diode D2 do not reflect
*physical devices but improve only modeling
*in the forward mode of operation.
*
.MODEL DIODE1 D
+ IS = 3E-16
+ N = 1.005
+ BV = {Vbreak}
+ IBV = 1E-09
+ RS = 0.05
+ CJO = 8.5E-11
+ VJ = 0.56
+ M = 0.324
+ FC = 0.5
+ TT = 0
+ EG = 1.1
+ XTI = 3
.MODEL DIODE2 D
+ IS = 7E-18
+ N = 1.25
+ RS = 8
.ENDS
*

